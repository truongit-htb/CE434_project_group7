`include "conv3d_kernel_3_channel_size_3.v"

module block1_conv1_8_kernel_3_channel #(
	parameter DATA_WIDTH = 32,
    parameter IMG_WIDTH = 56,
    parameter IMG_HEIGHT = 56,
    parameter SIZE = 3,
    parameter CHANNEL = 3,
    // parameter NUM_KERNEL = 8,

    // Kx_Cy_Wz = KERNELx_CHANNELy_WEIGHTz
    
	parameter K0_C0_W0 = 32'hbe5457b9,
	parameter K0_C0_W1 = 32'hbe550164,
	parameter K0_C0_W2 = 32'hbe2f75a6,
	parameter K0_C0_W3 = 32'hbe2f678b,
	parameter K0_C0_W4 = 32'hbe41dd65,
	parameter K0_C0_W5 = 32'hbe1cb911,
	parameter K0_C0_W6 = 32'h3e0f0fa3,
	parameter K0_C0_W7 = 32'h3e25c97c,
	parameter K0_C0_W8 = 32'h3d81a358,
	parameter K0_C1_W0 = 32'hbe55a967,
	parameter K0_C1_W1 = 32'hbd9429ce,
	parameter K0_C1_W2 = 32'h3c90fb11,
	parameter K0_C1_W3 = 32'h3dcbff4c,
	parameter K0_C1_W4 = 32'h3c90b7c4,
	parameter K0_C1_W5 = 32'h3e75047e,
	parameter K0_C1_W6 = 32'h3de8fd9e,
	parameter K0_C1_W7 = 32'h3e6056a7,
	parameter K0_C1_W8 = 32'h3e0a27e4,
	parameter K0_C2_W0 = 32'hbbb69696,
	parameter K0_C2_W1 = 32'h3e5f9c8c,
	parameter K0_C2_W2 = 32'hbe275eb2,
	parameter K0_C2_W3 = 32'hbdfb1afe,
	parameter K0_C2_W4 = 32'hbe66ea42,
	parameter K0_C2_W5 = 32'h3db88d53,
	parameter K0_C2_W6 = 32'hbccb4ca1,
	parameter K0_C2_W7 = 32'h3d9ff8a8,
	parameter K0_C2_W8 = 32'h3e2134bc,
	parameter K0_BIAS  = 32'h3ba40ddd,

	parameter K1_C0_W0 = 32'h3e6f7ea0,
	parameter K1_C0_W1 = 32'h3caea37a,
	parameter K1_C0_W2 = 32'h3e61a449,
	parameter K1_C0_W3 = 32'h3dfc7e86,
	parameter K1_C0_W4 = 32'h3e72c593,
	parameter K1_C0_W5 = 32'h3e40fdf8,
	parameter K1_C0_W6 = 32'h3d2b356f,
	parameter K1_C0_W7 = 32'hbd3d2302,
	parameter K1_C0_W8 = 32'hbdfd658e,
	parameter K1_C1_W0 = 32'hbd96d5e1,
	parameter K1_C1_W1 = 32'h3e49ad6b,
	parameter K1_C1_W2 = 32'hbe1c02c3,
	parameter K1_C1_W3 = 32'hbe275c3a,
	parameter K1_C1_W4 = 32'hbe6ccf39,
	parameter K1_C1_W5 = 32'h3e509fe9,
	parameter K1_C1_W6 = 32'hbe694c6a,
	parameter K1_C1_W7 = 32'hbd87850d,
	parameter K1_C1_W8 = 32'hbe250ae2,
	parameter K1_C2_W0 = 32'h3e369083,
	parameter K1_C2_W1 = 32'hbe4b95e0,
	parameter K1_C2_W2 = 32'h3df432cc,
	parameter K1_C2_W3 = 32'hbe05335a,
	parameter K1_C2_W4 = 32'h3e1f3ea7,
	parameter K1_C2_W5 = 32'hbe05a7a4,
	parameter K1_C2_W6 = 32'hbe30e846,
	parameter K1_C2_W7 = 32'h3e53f372,
	parameter K1_C2_W8 = 32'hbd88fe16,
	parameter K1_BIAS  = 32'hba54c9af,

	parameter K2_C0_W0 = 32'h3d07daba,
	parameter K2_C0_W1 = 32'hbe5c9335,
	parameter K2_C0_W2 = 32'h3e763928,
	parameter K2_C0_W3 = 32'hbe650b6c,
	parameter K2_C0_W4 = 32'h3e5d62ed,
	parameter K2_C0_W5 = 32'h3e049c9b,
	parameter K2_C0_W6 = 32'hbe395fb7,
	parameter K2_C0_W7 = 32'hbc0afd89,
	parameter K2_C0_W8 = 32'h3deacb0f,
	parameter K2_C1_W0 = 32'h3d9c27d8,
	parameter K2_C1_W1 = 32'h3e277674,
	parameter K2_C1_W2 = 32'h3daf8704,
	parameter K2_C1_W3 = 32'hbe0f9f2b,
	parameter K2_C1_W4 = 32'h397632dc,
	parameter K2_C1_W5 = 32'h3e672872,
	parameter K2_C1_W6 = 32'h3e6847bf,
	parameter K2_C1_W7 = 32'h3e4e17ba,
	parameter K2_C1_W8 = 32'hbe1ea955,
	parameter K2_C2_W0 = 32'hbe2d302d,
	parameter K2_C2_W1 = 32'hbe65988f,
	parameter K2_C2_W2 = 32'h3e67611e,
	parameter K2_C2_W3 = 32'hbe51c5b3,
	parameter K2_C2_W4 = 32'hbe60391b,
	parameter K2_C2_W5 = 32'hbe32e6e9,
	parameter K2_C2_W6 = 32'hbde2014e,
	parameter K2_C2_W7 = 32'h3cf93ae7,
	parameter K2_C2_W8 = 32'hbda29f21,
	parameter K2_BIAS  = 32'h3b4bd824,

	parameter K3_C0_W0 = 32'hbe52e23c,
	parameter K3_C0_W1 = 32'hbdeab053,
	parameter K3_C0_W2 = 32'hbe1b9e11,
	parameter K3_C0_W3 = 32'hbe0f264a,
	parameter K3_C0_W4 = 32'h3dc58431,
	parameter K3_C0_W5 = 32'h3e795a02,
	parameter K3_C0_W6 = 32'hbdddeaeb,
	parameter K3_C0_W7 = 32'h3e2bf964,
	parameter K3_C0_W8 = 32'h3e66cc48,
	parameter K3_C1_W0 = 32'hbdc2c8c6,
	parameter K3_C1_W1 = 32'hbdb3c262,
	parameter K3_C1_W2 = 32'h3e2006ea,
	parameter K3_C1_W3 = 32'h3d37c013,
	parameter K3_C1_W4 = 32'h3d3942d6,
	parameter K3_C1_W5 = 32'h3da2a61f,
	parameter K3_C1_W6 = 32'hbe6b533f,
	parameter K3_C1_W7 = 32'hbdd3ca4a,
	parameter K3_C1_W8 = 32'h3da37bbc,
	parameter K3_C2_W0 = 32'hbd996e27,
	parameter K3_C2_W1 = 32'h3e7187c4,
	parameter K3_C2_W2 = 32'hbe684669,
	parameter K3_C2_W3 = 32'h3d999772,
	parameter K3_C2_W4 = 32'h3c45466b,
	parameter K3_C2_W5 = 32'hbcfbb100,
	parameter K3_C2_W6 = 32'h3da09531,
	parameter K3_C2_W7 = 32'hbe3d3a62,
	parameter K3_C2_W8 = 32'h3d825f02,
	parameter K3_BIAS  = 32'h39541cad,

	parameter K4_C0_W0 = 32'hbe635d4a,
	parameter K4_C0_W1 = 32'hbe2d7633,
	parameter K4_C0_W2 = 32'hbd97f084,
	parameter K4_C0_W3 = 32'h3d17ff1a,
	parameter K4_C0_W4 = 32'hbda0c98c,
	parameter K4_C0_W5 = 32'hbcfd5a36,
	parameter K4_C0_W6 = 32'h3e523dc4,
	parameter K4_C0_W7 = 32'hbe399bfa,
	parameter K4_C0_W8 = 32'h3e57bdbb,
	parameter K4_C1_W0 = 32'hbd860e66,
	parameter K4_C1_W1 = 32'h3e344aac,
	parameter K4_C1_W2 = 32'h3e2a5bee,
	parameter K4_C1_W3 = 32'h3e23f378,
	parameter K4_C1_W4 = 32'hbdba45b1,
	parameter K4_C1_W5 = 32'h3de014f5,
	parameter K4_C1_W6 = 32'hbd1a1239,
	parameter K4_C1_W7 = 32'h3d5589f7,
	parameter K4_C1_W8 = 32'h3dffd925,
	parameter K4_C2_W0 = 32'h3d1f3a14,
	parameter K4_C2_W1 = 32'h3e73cdb0,
	parameter K4_C2_W2 = 32'hbe677a84,
	parameter K4_C2_W3 = 32'h3e4e7393,
	parameter K4_C2_W4 = 32'hbcf86179,
	parameter K4_C2_W5 = 32'h3dae562c,
	parameter K4_C2_W6 = 32'hbe0792e2,
	parameter K4_C2_W7 = 32'h3e68cee2,
	parameter K4_C2_W8 = 32'hbdbce6db,
	parameter K4_BIAS  = 32'h3a0c6cdb,

	parameter K5_C0_W0 = 32'hbe6cf90a,
	parameter K5_C0_W1 = 32'h3e5569a1,
	parameter K5_C0_W2 = 32'h3c5df7d5,
	parameter K5_C0_W3 = 32'h3da9607e,
	parameter K5_C0_W4 = 32'h3dcde027,
	parameter K5_C0_W5 = 32'h3e2538b2,
	parameter K5_C0_W6 = 32'hbd453418,
	parameter K5_C0_W7 = 32'h3e43c282,
	parameter K5_C0_W8 = 32'h3e2e2530,
	parameter K5_C1_W0 = 32'h3dacbfe7,
	parameter K5_C1_W1 = 32'h3e43263e,
	parameter K5_C1_W2 = 32'h3e20d66a,
	parameter K5_C1_W3 = 32'h3e048bbd,
	parameter K5_C1_W4 = 32'hbe69b4e6,
	parameter K5_C1_W5 = 32'h3e0d300b,
	parameter K5_C1_W6 = 32'h3df146f1,
	parameter K5_C1_W7 = 32'hbe66eabd,
	parameter K5_C1_W8 = 32'h3d64534e,
	parameter K5_C2_W0 = 32'hbe62f4a6,
	parameter K5_C2_W1 = 32'h3d839ee0,
	parameter K5_C2_W2 = 32'hbdb22566,
	parameter K5_C2_W3 = 32'h3d6d5dd5,
	parameter K5_C2_W4 = 32'hbe1977ac,
	parameter K5_C2_W5 = 32'hbdb233b1,
	parameter K5_C2_W6 = 32'h3e3915f0,
	parameter K5_C2_W7 = 32'hbe5c30fb,
	parameter K5_C2_W8 = 32'hbc0b443a,
	parameter K5_BIAS  = 32'hba88bac6,

	parameter K6_C0_W0 = 32'hbe4a448d,
	parameter K6_C0_W1 = 32'hbbe89ac5,
	parameter K6_C0_W2 = 32'hbd0eafd4,
	parameter K6_C0_W3 = 32'hbd4ef2d8,
	parameter K6_C0_W4 = 32'h3e452f0d,
	parameter K6_C0_W5 = 32'h3e20208e,
	parameter K6_C0_W6 = 32'h3d75d1d6,
	parameter K6_C0_W7 = 32'h3d4cbe78,
	parameter K6_C0_W8 = 32'hbde56c4d,
	parameter K6_C1_W0 = 32'h3e40e185,
	parameter K6_C1_W1 = 32'h3d295fe3,
	parameter K6_C1_W2 = 32'hbe32554e,
	parameter K6_C1_W3 = 32'h3e3d1005,
	parameter K6_C1_W4 = 32'h3d1d65d4,
	parameter K6_C1_W5 = 32'h3e734e38,
	parameter K6_C1_W6 = 32'hbd953dea,
	parameter K6_C1_W7 = 32'h3dd8ed00,
	parameter K6_C1_W8 = 32'h3e23aaa5,
	parameter K6_C2_W0 = 32'h3e53b7fa,
	parameter K6_C2_W1 = 32'h3df1e79b,
	parameter K6_C2_W2 = 32'h3e3da7f7,
	parameter K6_C2_W3 = 32'h3dcf6a7b,
	parameter K6_C2_W4 = 32'h3e1ff682,
	parameter K6_C2_W5 = 32'h3d3bb6ec,
	parameter K6_C2_W6 = 32'hbda45370,
	parameter K6_C2_W7 = 32'hbe33d8cf,
	parameter K6_C2_W8 = 32'h3df15b1d,
	parameter K6_BIAS  = 32'hbafbcb0c,

	parameter K7_C0_W0 = 32'h3e3c7e5d,
	parameter K7_C0_W1 = 32'h3d9228bd,
	parameter K7_C0_W2 = 32'hbe3bf8e7,
	parameter K7_C0_W3 = 32'h3d972aa7,
	parameter K7_C0_W4 = 32'hbe71610c,
	parameter K7_C0_W5 = 32'hbe1ecaa1,
	parameter K7_C0_W6 = 32'hbc6197ad,
	parameter K7_C0_W7 = 32'hbd185843,
	parameter K7_C0_W8 = 32'h3ccf49ee,
	parameter K7_C1_W0 = 32'hbe6bacf4,
	parameter K7_C1_W1 = 32'h3cb0ab15,
	parameter K7_C1_W2 = 32'h3e6d8037,
	parameter K7_C1_W3 = 32'hbd665558,
	parameter K7_C1_W4 = 32'h3e6080ac,
	parameter K7_C1_W5 = 32'hbe61b862,
	parameter K7_C1_W6 = 32'h3e331cda,
	parameter K7_C1_W7 = 32'hbe50cfb7,
	parameter K7_C1_W8 = 32'hbbf1a9e4,
	parameter K7_C2_W0 = 32'h3d8fa1ee,
	parameter K7_C2_W1 = 32'h3e1c5bf4,
	parameter K7_C2_W2 = 32'hbe79bebb,
	parameter K7_C2_W3 = 32'hbd6e4230,
	parameter K7_C2_W4 = 32'h3cb1ba57,
	parameter K7_C2_W5 = 32'hbe5831d8,
	parameter K7_C2_W6 = 32'h3e1f010d,
	parameter K7_C2_W7 = 32'h3d36a248,
	parameter K7_C2_W8 = 32'hbb56deb8,
	parameter K7_BIAS  = 32'h3bd0f0a8
    )
    (
    input     wire            clk,
    input     wire            resetn,
    input     wire            data_valid_in,
    input     wire   [DATA_WIDTH-1:0]    data_in0,
    input     wire   [DATA_WIDTH-1:0]    data_in1,
    input     wire   [DATA_WIDTH-1:0]    data_in2,
    
    output     wire   [DATA_WIDTH-1:0]    data_out_conv0,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv1,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv2,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv3,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv4,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv5,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv6,
    output     wire   [DATA_WIDTH-1:0]    data_out_conv7,

    output     valid_out_pixel,
    output reg done_img
    );

    reg [31:0] counter;
    wire valid_out_conv0, valid_out_conv1, valid_out_conv2, valid_out_conv3, valid_out_conv4, valid_out_conv5, valid_out_conv6, valid_out_conv7; 
	wire done_conv_0, done_conv_1, done_conv_2, done_conv_3, done_conv_4, done_conv_5, done_conv_6, done_conv_7; 

    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K0_C0_W0),
        .C0_W1(K0_C0_W1),
        .C0_W2(K0_C0_W2),
        .C0_W3(K0_C0_W3),
        .C0_W4(K0_C0_W4),
        .C0_W5(K0_C0_W5),
        .C0_W6(K0_C0_W6),
        .C0_W7(K0_C0_W7),
        .C0_W8(K0_C0_W8),
        .C1_W0(K0_C1_W0),
        .C1_W1(K0_C1_W1),
        .C1_W2(K0_C1_W2),
        .C1_W3(K0_C1_W3),
        .C1_W4(K0_C1_W4),
        .C1_W5(K0_C1_W5),
        .C1_W6(K0_C1_W6),
        .C1_W7(K0_C1_W7),
        .C1_W8(K0_C1_W8),
        .C2_W0(K0_C2_W0),
        .C2_W1(K0_C2_W1),
        .C2_W2(K0_C2_W2),
        .C2_W3(K0_C2_W3),
        .C2_W4(K0_C2_W4),
        .C2_W5(K0_C2_W5),
        .C2_W6(K0_C2_W6),
        .C2_W7(K0_C2_W7),
        .C2_W8(K0_C2_W8),
        .BIAS(K0_BIAS)
		)
		conv1_0(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,            
		data_out_conv0,
		valid_out_conv0,
		done_conv_0
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K1_C0_W0),
        .C0_W1(K1_C0_W1),
        .C0_W2(K1_C0_W2),
        .C0_W3(K1_C0_W3),
        .C0_W4(K1_C0_W4),
        .C0_W5(K1_C0_W5),
        .C0_W6(K1_C0_W6),
        .C0_W7(K1_C0_W7),
        .C0_W8(K1_C0_W8),
        .C1_W0(K1_C1_W0),
        .C1_W1(K1_C1_W1),
        .C1_W2(K1_C1_W2),
        .C1_W3(K1_C1_W3),
        .C1_W4(K1_C1_W4),
        .C1_W5(K1_C1_W5),
        .C1_W6(K1_C1_W6),
        .C1_W7(K1_C1_W7),
        .C1_W8(K1_C1_W8),
        .C2_W0(K1_C2_W0),
        .C2_W1(K1_C2_W1),
        .C2_W2(K1_C2_W2),
        .C2_W3(K1_C2_W3),
        .C2_W4(K1_C2_W4),
        .C2_W5(K1_C2_W5),
        .C2_W6(K1_C2_W6),
        .C2_W7(K1_C2_W7),
        .C2_W8(K1_C2_W8),
        .BIAS(K1_BIAS)
		)
		conv1_1(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,   
		data_out_conv1,
		valid_out_conv1,
		done_conv_1
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K2_C0_W0),
        .C0_W1(K2_C0_W1),
        .C0_W2(K2_C0_W2),
        .C0_W3(K2_C0_W3),
        .C0_W4(K2_C0_W4),
        .C0_W5(K2_C0_W5),
        .C0_W6(K2_C0_W6),
        .C0_W7(K2_C0_W7),
        .C0_W8(K2_C0_W8),
        .C1_W0(K2_C1_W0),
        .C1_W1(K2_C1_W1),
        .C1_W2(K2_C1_W2),
        .C1_W3(K2_C1_W3),
        .C1_W4(K2_C1_W4),
        .C1_W5(K2_C1_W5),
        .C1_W6(K2_C1_W6),
        .C1_W7(K2_C1_W7),
        .C1_W8(K2_C1_W8),
        .C2_W0(K2_C2_W0),
        .C2_W1(K2_C2_W1),
        .C2_W2(K2_C2_W2),
        .C2_W3(K2_C2_W3),
        .C2_W4(K2_C2_W4),
        .C2_W5(K2_C2_W5),
        .C2_W6(K2_C2_W6),
        .C2_W7(K2_C2_W7),
        .C2_W8(K2_C2_W8),
        .BIAS(K2_BIAS)
		)
		conv1_2(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,   
		data_out_conv2,
		valid_out_conv2,
		done_conv_2
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K3_C0_W0),
        .C0_W1(K3_C0_W1),
        .C0_W2(K3_C0_W2),
        .C0_W3(K3_C0_W3),
        .C0_W4(K3_C0_W4),
        .C0_W5(K3_C0_W5),
        .C0_W6(K3_C0_W6),
        .C0_W7(K3_C0_W7),
        .C0_W8(K3_C0_W8),
        .C1_W0(K3_C1_W0),
        .C1_W1(K3_C1_W1),
        .C1_W2(K3_C1_W2),
        .C1_W3(K3_C1_W3),
        .C1_W4(K3_C1_W4),
        .C1_W5(K3_C1_W5),
        .C1_W6(K3_C1_W6),
        .C1_W7(K3_C1_W7),
        .C1_W8(K3_C1_W8),
        .C2_W0(K3_C2_W0),
        .C2_W1(K3_C2_W1),
        .C2_W2(K3_C2_W2),
        .C2_W3(K3_C2_W3),
        .C2_W4(K3_C2_W4),
        .C2_W5(K3_C2_W5),
        .C2_W6(K3_C2_W6),
        .C2_W7(K3_C2_W7),
        .C2_W8(K3_C2_W8),
        .BIAS(K3_BIAS)
		)
		conv1_3(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,
		data_out_conv3,
		valid_out_conv3,
		done_conv_3
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K4_C0_W0),
        .C0_W1(K4_C0_W1),
        .C0_W2(K4_C0_W2),
        .C0_W3(K4_C0_W3),
        .C0_W4(K4_C0_W4),
        .C0_W5(K4_C0_W5),
        .C0_W6(K4_C0_W6),
        .C0_W7(K4_C0_W7),
        .C0_W8(K4_C0_W8),
        .C1_W0(K4_C1_W0),
        .C1_W1(K4_C1_W1),
        .C1_W2(K4_C1_W2),
        .C1_W3(K4_C1_W3),
        .C1_W4(K4_C1_W4),
        .C1_W5(K4_C1_W5),
        .C1_W6(K4_C1_W6),
        .C1_W7(K4_C1_W7),
        .C1_W8(K4_C1_W8),
        .C2_W0(K4_C2_W0),
        .C2_W1(K4_C2_W1),
        .C2_W2(K4_C2_W2),
        .C2_W3(K4_C2_W3),
        .C2_W4(K4_C2_W4),
        .C2_W5(K4_C2_W5),
        .C2_W6(K4_C2_W6),
        .C2_W7(K4_C2_W7),
        .C2_W8(K4_C2_W8),
        .BIAS(K4_BIAS)
		)
		conv1_4(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,  
		data_out_conv4,
		valid_out_conv4,
		done_conv_4
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K5_C0_W0),
        .C0_W1(K5_C0_W1),
        .C0_W2(K5_C0_W2),
        .C0_W3(K5_C0_W3),
        .C0_W4(K5_C0_W4),
        .C0_W5(K5_C0_W5),
        .C0_W6(K5_C0_W6),
        .C0_W7(K5_C0_W7),
        .C0_W8(K5_C0_W8),
        .C1_W0(K5_C1_W0),
        .C1_W1(K5_C1_W1),
        .C1_W2(K5_C1_W2),
        .C1_W3(K5_C1_W3),
        .C1_W4(K5_C1_W4),
        .C1_W5(K5_C1_W5),
        .C1_W6(K5_C1_W6),
        .C1_W7(K5_C1_W7),
        .C1_W8(K5_C1_W8),
        .C2_W0(K5_C2_W0),
        .C2_W1(K5_C2_W1),
        .C2_W2(K5_C2_W2),
        .C2_W3(K5_C2_W3),
        .C2_W4(K5_C2_W4),
        .C2_W5(K5_C2_W5),
        .C2_W6(K5_C2_W6),
        .C2_W7(K5_C2_W7),
        .C2_W8(K5_C2_W8),
        .BIAS(K5_BIAS)
		)
		conv1_5(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,        
		data_out_conv5,
		valid_out_conv5,
		done_conv_5
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K6_C0_W0),
        .C0_W1(K6_C0_W1),
        .C0_W2(K6_C0_W2),
        .C0_W3(K6_C0_W3),
        .C0_W4(K6_C0_W4),
        .C0_W5(K6_C0_W5),
        .C0_W6(K6_C0_W6),
        .C0_W7(K6_C0_W7),
        .C0_W8(K6_C0_W8),
        .C1_W0(K6_C1_W0),
        .C1_W1(K6_C1_W1),
        .C1_W2(K6_C1_W2),
        .C1_W3(K6_C1_W3),
        .C1_W4(K6_C1_W4),
        .C1_W5(K6_C1_W5),
        .C1_W6(K6_C1_W6),
        .C1_W7(K6_C1_W7),
        .C1_W8(K6_C1_W8),
        .C2_W0(K6_C2_W0),
        .C2_W1(K6_C2_W1),
        .C2_W2(K6_C2_W2),
        .C2_W3(K6_C2_W3),
        .C2_W4(K6_C2_W4),
        .C2_W5(K6_C2_W5),
        .C2_W6(K6_C2_W6),
        .C2_W7(K6_C2_W7),
        .C2_W8(K6_C2_W8),
        .BIAS(K6_BIAS)
		)
		conv1_6(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,
		data_out_conv6,
		valid_out_conv6,
		done_conv_6
		);
    conv3d_kernel_3_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(IMG_WIDTH),.IMG_HEIGHT(IMG_HEIGHT),
        .C0_W0(K7_C0_W0),
        .C0_W1(K7_C0_W1),
        .C0_W2(K7_C0_W2),
        .C0_W3(K7_C0_W3),
        .C0_W4(K7_C0_W4),
        .C0_W5(K7_C0_W5),
        .C0_W6(K7_C0_W6),
        .C0_W7(K7_C0_W7),
        .C0_W8(K7_C0_W8),
        .C1_W0(K7_C1_W0),
        .C1_W1(K7_C1_W1),
        .C1_W2(K7_C1_W2),
        .C1_W3(K7_C1_W3),
        .C1_W4(K7_C1_W4),
        .C1_W5(K7_C1_W5),
        .C1_W6(K7_C1_W6),
        .C1_W7(K7_C1_W7),
        .C1_W8(K7_C1_W8),
        .C2_W0(K7_C2_W0),
        .C2_W1(K7_C2_W1),
        .C2_W2(K7_C2_W2),
        .C2_W3(K7_C2_W3),
        .C2_W4(K7_C2_W4),
        .C2_W5(K7_C2_W5),
        .C2_W6(K7_C2_W6),
        .C2_W7(K7_C2_W7),
        .C2_W8(K7_C2_W8),
        .BIAS(K7_BIAS)
		)
		conv1_7(
		clk,
		resetn,
		data_valid_in,
		data_in0,
        data_in1,
        data_in2,    
		data_out_conv7,
		valid_out_conv7,
		done_conv_7
		);

    assign valid_out_pixel = valid_out_conv7;
    
    always @ (posedge clk or negedge resetn) 
    begin
        if(resetn == 1'b0) 
            counter <= 0;
        else 
            if (done_img == 1'b1) begin
                counter <= 0;
            end
            else 
                if(valid_out_pixel == 1'b1) 
                begin
                    if(counter == (IMG_WIDTH)*(IMG_HEIGHT) -1 ) 
                        counter <= 0;
                    else 
                        counter <= counter + 1;
                end
                else 
                    counter <= counter;
    end

    always @ (posedge clk or negedge resetn) 
    begin
        if(resetn == 1'b0) 
            done_img <= 0;
        else 
            if(counter == (IMG_WIDTH)*(IMG_HEIGHT) -2) 
                done_img <= (valid_out_pixel)?1'b1:1'b0;
            else 
                done_img <= 0;
    end

endmodule