`ifndef ACTIVATE_INCLUDED
    `include "activate.v"
    `define ACTIVATE_INCLUDED
`endif
`ifndef MAX_POOLING_INCLUDED
    `include "max_pooling.v"
    `define MAX_POOLING_INCLUDED
`endif

module block_demo #(
    parameter DATA_WIDTH = 32,
    parameter WIDTH = 56,
    parameter HEIGHT = 56,
    parameter CHANNEL_OUT = 16
    ) 
    (
    input	clk,
	input	resetn,
	input	valid_in,
	input	[DATA_WIDTH-1:0]	data_in_0,
	input	[DATA_WIDTH-1:0]	data_in_1,
	input	[DATA_WIDTH-1:0]	data_in_2,
	input	[DATA_WIDTH-1:0]	data_in_3,
	input	[DATA_WIDTH-1:0]	data_in_4,
	input	[DATA_WIDTH-1:0]	data_in_5,
	input	[DATA_WIDTH-1:0]	data_in_6,
	input	[DATA_WIDTH-1:0]	data_in_7,
	output	[DATA_WIDTH-1:0]	data_out_0,
	output	[DATA_WIDTH-1:0]	data_out_1,
	output	[DATA_WIDTH-1:0]	data_out_2,
	output	[DATA_WIDTH-1:0]	data_out_3,
	output	[DATA_WIDTH-1:0]	data_out_4,
	output	[DATA_WIDTH-1:0]	data_out_5,
	output	[DATA_WIDTH-1:0]	data_out_6,
	output	[DATA_WIDTH-1:0]	data_out_7,
	output	[DATA_WIDTH-1:0]	data_out_8,
	output	[DATA_WIDTH-1:0]	data_out_9,
	output	[DATA_WIDTH-1:0]	data_out_10,
	output	[DATA_WIDTH-1:0]	data_out_11,
	output	[DATA_WIDTH-1:0]	data_out_12,
	output	[DATA_WIDTH-1:0]	data_out_13,
	output	[DATA_WIDTH-1:0]	data_out_14,
	output	[DATA_WIDTH-1:0]	data_out_15,
	output	valid_out,
	output	done
    );

    wire [DATA_WIDTH-1:0] conv_out_4_1  [0: CHANNEL_OUT -1];    
    wire conv_valid_out_4_1;
    wire done_conv_4_1;

    wire [DATA_WIDTH-1:0] conv_out_4_2  [0: CHANNEL_OUT -1];    
    wire conv_valid_out_4_2;
    wire done_conv_4_2;

	wire [DATA_WIDTH-1:0] conv_out_4_3  [0: CHANNEL_OUT -1];    
    wire conv_valid_out_4_3;
    wire done_conv_4_3;


    // WITH RELU AND MAX_POOLING
    wire [DATA_WIDTH-1:0] relu_out  [0: CHANNEL_OUT -1];

    wire [DATA_WIDTH-1:0] data_out_pool [0: CHANNEL_OUT -1];
    wire [CHANNEL_OUT -1 : 0] valid_out_pool;
    wire [CHANNEL_OUT -1 : 0] done_pool;
    
    assign data_out_0 = data_out_pool[0];
    assign data_out_1 = data_out_pool[1];
    assign data_out_2 = data_out_pool[2];
    assign data_out_3 = data_out_pool[3];
    assign data_out_4 = data_out_pool[4];
    assign data_out_5 = data_out_pool[5];
    assign data_out_6 = data_out_pool[6];
    assign data_out_7 = data_out_pool[7];
    assign data_out_8 = data_out_pool[8];
	assign data_out_9 = data_out_pool[9];
	assign data_out_10 = data_out_pool[10];
	assign data_out_11 = data_out_pool[11];
	assign data_out_12 = data_out_pool[12];
	assign data_out_13 = data_out_pool[13];
	assign data_out_14 = data_out_pool[14];
	assign data_out_15 = data_out_pool[15];

    assign valid_out = valid_out_pool[CHANNEL_OUT -1];
    assign done = done_pool[CHANNEL_OUT -1];
    // -------------------------------------



    // ONLY CONV - WITHOUT RELU AND MAX_POOLING
    // assign valid_out = conv_valid_out_4_2;	// Edit here
    // assign done = done_conv_4_2;				// Edit here

    // assign data_out_0 = conv_out_4_2[0];
	// assign data_out_1 = conv_out_4_2[1];
	// assign data_out_2 = conv_out_4_2[2];
	// assign data_out_3 = conv_out_4_2[3];
	// assign data_out_4 = conv_out_4_2[4];
	// assign data_out_5 = conv_out_4_2[5];
	// assign data_out_6 = conv_out_4_2[6];
	// assign data_out_7 = conv_out_4_2[7];
	// assign data_out_8 = conv_out_4_2[8];
	// assign data_out_9 = conv_out_4_2[9];
	// assign data_out_10 = conv_out_4_2[10];
	// assign data_out_11 = conv_out_4_2[11];
	// assign data_out_12 = conv_out_4_2[12];
	// assign data_out_13 = conv_out_4_2[13];
	// assign data_out_14 = conv_out_4_2[14];
	// assign data_out_15 = conv_out_4_2[15];
    // -------------------------------------


	conv3d_16_kernel_8_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(WIDTH),.IMG_HEIGHT(HEIGHT),
		.K0_C0_W0(32'h3d3f35fd), .K0_C0_W1(32'h3d811f77), .K0_C0_W2(32'hbe1d022a), .K0_C0_W3(32'h3e161386), .K0_C0_W4(32'h3d1a89c4), .K0_C0_W5(32'h3db4d8a3), .K0_C0_W6(32'h3e0e3a1a), .K0_C0_W7(32'h3cc9dd22), .K0_C0_W8(32'hbe34e767), 
		.K0_C1_W0(32'hbcbbcb57), .K0_C1_W1(32'h3dae3dca), .K0_C1_W2(32'h3c905611), .K0_C1_W3(32'hbc847bed), .K0_C1_W4(32'hbd61f3a6), .K0_C1_W5(32'hbda9bab2), .K0_C1_W6(32'hbd45a29e), .K0_C1_W7(32'hbe31d201), .K0_C1_W8(32'h3d79d165), 
		.K0_C2_W0(32'h3e5b6f5b), .K0_C2_W1(32'h3d253094), .K0_C2_W2(32'hbda1a404), .K0_C2_W3(32'h3d8586f9), .K0_C2_W4(32'hbd07c599), .K0_C2_W5(32'h3dfb1b50), .K0_C2_W6(32'h3dbb036d), .K0_C2_W7(32'hbdc29740), .K0_C2_W8(32'h3d214c8c), 
		.K0_C3_W0(32'h3e447eae), .K0_C3_W1(32'hbd3bb6d5), .K0_C3_W2(32'h3d8dd03f), .K0_C3_W3(32'hbd8f6fc4), .K0_C3_W4(32'h3da6db66), .K0_C3_W5(32'h3dd33b70), .K0_C3_W6(32'h3e26c7e7), .K0_C3_W7(32'h3df61a28), .K0_C3_W8(32'h3d84f053), 
		.K0_C4_W0(32'h3e325a9e), .K0_C4_W1(32'h3d8c3135), .K0_C4_W2(32'h3d963617), .K0_C4_W3(32'hbb683e92), .K0_C4_W4(32'h3cdef154), .K0_C4_W5(32'h3dc4b775), .K0_C4_W6(32'hbd1b4cab), .K0_C4_W7(32'h3d8cdf3e), .K0_C4_W8(32'h3e00bc05), 
		.K0_C5_W0(32'h3e12961a), .K0_C5_W1(32'hbdd01ec4), .K0_C5_W2(32'hbcc46adf), .K0_C5_W3(32'h3c8d2e91), .K0_C5_W4(32'hbe4222b9), .K0_C5_W5(32'hbd55e588), .K0_C5_W6(32'h3d501afd), .K0_C5_W7(32'hbe2271fd), .K0_C5_W8(32'hbe1958fc), 
		.K0_C6_W0(32'hbe0ea4a4), .K0_C6_W1(32'hbd3a00ca), .K0_C6_W2(32'h3e0d752c), .K0_C6_W3(32'hbe20584c), .K0_C6_W4(32'h3db49aec), .K0_C6_W5(32'h3d1ab6fd), .K0_C6_W6(32'hbdc2c87d), .K0_C6_W7(32'h3e2310aa), .K0_C6_W8(32'hbda25e0b), 
		.K0_C7_W0(32'h3d2dfc15), .K0_C7_W1(32'h3e04f176), .K0_C7_W2(32'h3daaa9b4), .K0_C7_W3(32'h3dfc30ef), .K0_C7_W4(32'hbd1da773), .K0_C7_W5(32'hbdf3e429), .K0_C7_W6(32'hbdfc99e3), .K0_C7_W7(32'hbe2c8330), .K0_C7_W8(32'hbe228cdf), 
		.K0_BIAS (32'hbd2963c5),

		.K1_C0_W0(32'h3bf5f6e0), .K1_C0_W1(32'h3dc4b5ba), .K1_C0_W2(32'hbd464263), .K1_C0_W3(32'h3dceb546), .K1_C0_W4(32'hbd968c86), .K1_C0_W5(32'hbb9ae053), .K1_C0_W6(32'hbe0185ee), .K1_C0_W7(32'hbdac3667), .K1_C0_W8(32'hbd22cba5), 
		.K1_C1_W0(32'h3b7a25b1), .K1_C1_W1(32'h3e41d0b9), .K1_C1_W2(32'hbd6a762c), .K1_C1_W3(32'hbc8d6d2b), .K1_C1_W4(32'hbcf35a5c), .K1_C1_W5(32'hbd2ca837), .K1_C1_W6(32'h3e3798a2), .K1_C1_W7(32'h3df673b4), .K1_C1_W8(32'h3d00648f), 
		.K1_C2_W0(32'hbe16525c), .K1_C2_W1(32'hbe0d14dd), .K1_C2_W2(32'h3d72954d), .K1_C2_W3(32'hbe058c7d), .K1_C2_W4(32'hbe40f228), .K1_C2_W5(32'hbdcff9f7), .K1_C2_W6(32'hbd386cd6), .K1_C2_W7(32'hbbae557d), .K1_C2_W8(32'h3b67c301), 
		.K1_C3_W0(32'h3dcadaf5), .K1_C3_W1(32'hbd48409b), .K1_C3_W2(32'hbc3e2551), .K1_C3_W3(32'hbb93be82), .K1_C3_W4(32'hbe0cff6c), .K1_C3_W5(32'hbdeaf903), .K1_C3_W6(32'hbd8664bc), .K1_C3_W7(32'hbd2ad5ca), .K1_C3_W8(32'h3d95dd5c), 
		.K1_C4_W0(32'hbcb7bcc3), .K1_C4_W1(32'h3cc586e0), .K1_C4_W2(32'h3dba60b5), .K1_C4_W3(32'h3db93869), .K1_C4_W4(32'h3cdbd72e), .K1_C4_W5(32'h3cb08afb), .K1_C4_W6(32'hbd7172bd), .K1_C4_W7(32'hbdba50a3), .K1_C4_W8(32'hbd1389e9), 
		.K1_C5_W0(32'h3c8b98fb), .K1_C5_W1(32'h3e36fee3), .K1_C5_W2(32'h3dc51262), .K1_C5_W3(32'hbdaa8a3b), .K1_C5_W4(32'h3e5a0217), .K1_C5_W5(32'hbe1e3695), .K1_C5_W6(32'hbd16faf3), .K1_C5_W7(32'hbce0e489), .K1_C5_W8(32'hbe02ba37), 
		.K1_C6_W0(32'hbe1adca8), .K1_C6_W1(32'hbd80871e), .K1_C6_W2(32'h3dce5259), .K1_C6_W3(32'h3d3a7da3), .K1_C6_W4(32'hbcbf8fe1), .K1_C6_W5(32'hbe087476), .K1_C6_W6(32'hbdaae47c), .K1_C6_W7(32'h3e1c1a64), .K1_C6_W8(32'hbc284315), 
		.K1_C7_W0(32'h3d9c4b00), .K1_C7_W1(32'hbd6d6edc), .K1_C7_W2(32'hbda8efc8), .K1_C7_W3(32'h3db060ae), .K1_C7_W4(32'h3b045649), .K1_C7_W5(32'hbe25fc5f), .K1_C7_W6(32'h3d0dc39d), .K1_C7_W7(32'hbd85d5ac), .K1_C7_W8(32'hbcb05310), 
		.K1_BIAS (32'h3d04c919),

		.K2_C0_W0(32'hbca95003), .K2_C0_W1(32'hbdaaa070), .K2_C0_W2(32'h3e0aeeb5), .K2_C0_W3(32'h3b085408), .K2_C0_W4(32'hbd926adc), .K2_C0_W5(32'hbdabdf09), .K2_C0_W6(32'h3df13ebb), .K2_C0_W7(32'hbd4e75f0), .K2_C0_W8(32'hbdc23856), 
		.K2_C1_W0(32'hbd472d12), .K2_C1_W1(32'hbdf98b7e), .K2_C1_W2(32'h3e27dc35), .K2_C1_W3(32'h3d64ff4e), .K2_C1_W4(32'h3c2dd180), .K2_C1_W5(32'h3e30d316), .K2_C1_W6(32'hbdddb8c0), .K2_C1_W7(32'h3e03dd7d), .K2_C1_W8(32'hbd9bec0a), 
		.K2_C2_W0(32'hbdbee88b), .K2_C2_W1(32'hbd31bf9b), .K2_C2_W2(32'hbdf143d2), .K2_C2_W3(32'hbdd4acb1), .K2_C2_W4(32'h3dfe1706), .K2_C2_W5(32'h3e3af9cc), .K2_C2_W6(32'h3d090965), .K2_C2_W7(32'hbe114c48), .K2_C2_W8(32'hbe213dfb), 
		.K2_C3_W0(32'hbae15dda), .K2_C3_W1(32'hbe17b4b7), .K2_C3_W2(32'hbe32f31d), .K2_C3_W3(32'h3d9312cc), .K2_C3_W4(32'h3b72f034), .K2_C3_W5(32'h3d96eb02), .K2_C3_W6(32'hbd5bc10b), .K2_C3_W7(32'hbe1221f1), .K2_C3_W8(32'h3d829cdb), 
		.K2_C4_W0(32'hbdbe68a5), .K2_C4_W1(32'hbe16ab93), .K2_C4_W2(32'h3e088fd7), .K2_C4_W3(32'h3cb1ebcd), .K2_C4_W4(32'hbcaed313), .K2_C4_W5(32'hbded3f19), .K2_C4_W6(32'hbdc3bea4), .K2_C4_W7(32'hbcdbeea4), .K2_C4_W8(32'hbe02392c), 
		.K2_C5_W0(32'hbddebc72), .K2_C5_W1(32'h3d6c6eeb), .K2_C5_W2(32'hbdf37409), .K2_C5_W3(32'h3deb3256), .K2_C5_W4(32'h3cbb7b7e), .K2_C5_W5(32'h3e1248e2), .K2_C5_W6(32'h3db98d79), .K2_C5_W7(32'hbe25699a), .K2_C5_W8(32'hbe10fb49), 
		.K2_C6_W0(32'h3d8783a8), .K2_C6_W1(32'h3d235240), .K2_C6_W2(32'h3d3fafd1), .K2_C6_W3(32'hbe12e773), .K2_C6_W4(32'hbd5b7fb9), .K2_C6_W5(32'hbdb933b6), .K2_C6_W6(32'hbdc976f9), .K2_C6_W7(32'h3df74e05), .K2_C6_W8(32'h3e24f268), 
		.K2_C7_W0(32'hbe25e90b), .K2_C7_W1(32'hbe24087d), .K2_C7_W2(32'h3d89a449), .K2_C7_W3(32'hbe0d6682), .K2_C7_W4(32'h3e120168), .K2_C7_W5(32'h3dfd1c5c), .K2_C7_W6(32'hbd096230), .K2_C7_W7(32'hbdd01420), .K2_C7_W8(32'h3d7528b1), 
		.K2_BIAS (32'h3d4b2c00),

		.K3_C0_W0(32'h3c2c4231), .K3_C0_W1(32'h3dec1be4), .K3_C0_W2(32'h3e5a8eed), .K3_C0_W3(32'hbe1c1a30), .K3_C0_W4(32'hbddb2cd5), .K3_C0_W5(32'h3dbd2fe0), .K3_C0_W6(32'hbd3e1e51), .K3_C0_W7(32'hbd932813), .K3_C0_W8(32'hbe2baeab), 
		.K3_C1_W0(32'h3d9658ba), .K3_C1_W1(32'hbc6380d5), .K3_C1_W2(32'h3db2100e), .K3_C1_W3(32'hbc8210d6), .K3_C1_W4(32'hbd9a2fc4), .K3_C1_W5(32'h3c0eae2c), .K3_C1_W6(32'hbd861ab4), .K3_C1_W7(32'h3dad79d7), .K3_C1_W8(32'h3ced611b), 
		.K3_C2_W0(32'hbd5092bb), .K3_C2_W1(32'h3d0a3132), .K3_C2_W2(32'h3db03663), .K3_C2_W3(32'hbda3f5e9), .K3_C2_W4(32'hbdba9faf), .K3_C2_W5(32'hbe1878f1), .K3_C2_W6(32'hbc8c2be4), .K3_C2_W7(32'h3c2dbdc5), .K3_C2_W8(32'h3cd46a28), 
		.K3_C3_W0(32'hbd8c5cf2), .K3_C3_W1(32'hbe331ce4), .K3_C3_W2(32'hbd596579), .K3_C3_W3(32'h3d82abb1), .K3_C3_W4(32'h3deac40f), .K3_C3_W5(32'h3e0bafef), .K3_C3_W6(32'hbe30690d), .K3_C3_W7(32'hbd764d36), .K3_C3_W8(32'hbdacc4c2), 
		.K3_C4_W0(32'hbe1843ac), .K3_C4_W1(32'h3dd32cff), .K3_C4_W2(32'hbe0441cf), .K3_C4_W3(32'h3c9ea3ea), .K3_C4_W4(32'h3d0930ef), .K3_C4_W5(32'h3c824841), .K3_C4_W6(32'h3e0b1df4), .K3_C4_W7(32'hbdb72356), .K3_C4_W8(32'h3da97b9c), 
		.K3_C5_W0(32'hbde69efe), .K3_C5_W1(32'hbd76959b), .K3_C5_W2(32'h3d0d43cb), .K3_C5_W3(32'h3e0641e7), .K3_C5_W4(32'hbd264aa1), .K3_C5_W5(32'hbc2f186b), .K3_C5_W6(32'h3e25afe7), .K3_C5_W7(32'h3d08bfc4), .K3_C5_W8(32'h3d34b8af), 
		.K3_C6_W0(32'h3d56e21c), .K3_C6_W1(32'hbdb74610), .K3_C6_W2(32'hbe2a12c6), .K3_C6_W3(32'h3e12c031), .K3_C6_W4(32'h3d8d1d97), .K3_C6_W5(32'h3de375f9), .K3_C6_W6(32'hbe46e08c), .K3_C6_W7(32'hbe3f5073), .K3_C6_W8(32'hbe0d6948), 
		.K3_C7_W0(32'h3e426426), .K3_C7_W1(32'h3cddc4ab), .K3_C7_W2(32'hbd8029d4), .K3_C7_W3(32'h3d75a2f8), .K3_C7_W4(32'hbd8040e2), .K3_C7_W5(32'hbe06d189), .K3_C7_W6(32'hbe126bd4), .K3_C7_W7(32'hbcf76c11), .K3_C7_W8(32'h3d79c02b), 
		.K3_BIAS (32'h3c5148c7),

		.K4_C0_W0(32'h3df1f6f2), .K4_C0_W1(32'hbdd37c65), .K4_C0_W2(32'hbe236573), .K4_C0_W3(32'h3ca965ca), .K4_C0_W4(32'h3e17ec14), .K4_C0_W5(32'h3e1555ff), .K4_C0_W6(32'h3e155505), .K4_C0_W7(32'hbdab320b), .K4_C0_W8(32'hbdfeeaa3), 
		.K4_C1_W0(32'h3cf9ff82), .K4_C1_W1(32'h3da38e9e), .K4_C1_W2(32'h3d82a660), .K4_C1_W3(32'h3d87b79c), .K4_C1_W4(32'hbd72b386), .K4_C1_W5(32'h3c7b95a8), .K4_C1_W6(32'h3e07b5b1), .K4_C1_W7(32'h3e050319), .K4_C1_W8(32'h3d56b4e0), 
		.K4_C2_W0(32'hbc527012), .K4_C2_W1(32'h3aa0626d), .K4_C2_W2(32'h3cd6259b), .K4_C2_W3(32'h3c8fa69d), .K4_C2_W4(32'hbd8c9751), .K4_C2_W5(32'h3d15d4f5), .K4_C2_W6(32'h3dcc8c96), .K4_C2_W7(32'h3d92783b), .K4_C2_W8(32'h3d2f1be2), 
		.K4_C3_W0(32'h3d152b7f), .K4_C3_W1(32'h3c6db8e0), .K4_C3_W2(32'hbd1170db), .K4_C3_W3(32'h3dc6eaa5), .K4_C3_W4(32'hbddbac56), .K4_C3_W5(32'h3d267892), .K4_C3_W6(32'h3dbca7fb), .K4_C3_W7(32'h3e2265d8), .K4_C3_W8(32'h3e0d1342), 
		.K4_C4_W0(32'hbdb6b787), .K4_C4_W1(32'h3d4171e3), .K4_C4_W2(32'hbbe23058), .K4_C4_W3(32'hbdb8905c), .K4_C4_W4(32'h3d838382), .K4_C4_W5(32'hbb39ca0a), .K4_C4_W6(32'h3c249639), .K4_C4_W7(32'h3dc9f974), .K4_C4_W8(32'h3d62b9c7), 
		.K4_C5_W0(32'hbd07d229), .K4_C5_W1(32'hbc3353bd), .K4_C5_W2(32'hbd932e43), .K4_C5_W3(32'hbe16a328), .K4_C5_W4(32'h3e02707e), .K4_C5_W5(32'hbd7387eb), .K4_C5_W6(32'hbc2399d5), .K4_C5_W7(32'h3d65b6b3), .K4_C5_W8(32'hbcf7be7c), 
		.K4_C6_W0(32'hbdc98b64), .K4_C6_W1(32'h3e27d45a), .K4_C6_W2(32'hbdcbda86), .K4_C6_W3(32'hbdd1c454), .K4_C6_W4(32'hbdefa5ec), .K4_C6_W5(32'h3dcd947a), .K4_C6_W6(32'hbe0791a8), .K4_C6_W7(32'hbe05c53c), .K4_C6_W8(32'hbcb4d981), 
		.K4_C7_W0(32'h3df5ecc8), .K4_C7_W1(32'hbd79ac62), .K4_C7_W2(32'h3e20a1b9), .K4_C7_W3(32'h3cac2d29), .K4_C7_W4(32'h3c7c36d1), .K4_C7_W5(32'hbd8a3a46), .K4_C7_W6(32'hbd45804b), .K4_C7_W7(32'hbe101264), .K4_C7_W8(32'h3dbe7d12), 
		.K4_BIAS (32'hbd85273a),

		.K5_C0_W0(32'hbdbf24d9), .K5_C0_W1(32'hbe1c860b), .K5_C0_W2(32'h3cf77d2f), .K5_C0_W3(32'h3e2b095a), .K5_C0_W4(32'h3db6145d), .K5_C0_W5(32'hbe2fe021), .K5_C0_W6(32'h3d5ae3eb), .K5_C0_W7(32'hbdf2ff18), .K5_C0_W8(32'h3d5944a4), 
		.K5_C1_W0(32'h3d4c42b2), .K5_C1_W1(32'h3df90696), .K5_C1_W2(32'hbd856212), .K5_C1_W3(32'h3dcbf3f7), .K5_C1_W4(32'h3e36bb6b), .K5_C1_W5(32'hbdfbd6ad), .K5_C1_W6(32'h3c6a7bfc), .K5_C1_W7(32'h3dfef6c2), .K5_C1_W8(32'h3da27fc2), 
		.K5_C2_W0(32'h3d156aa9), .K5_C2_W1(32'hbc168d5b), .K5_C2_W2(32'hbd93504e), .K5_C2_W3(32'hbd047d99), .K5_C2_W4(32'h3d5f4028), .K5_C2_W5(32'hbe448ceb), .K5_C2_W6(32'hbd9a7e09), .K5_C2_W7(32'hbe483566), .K5_C2_W8(32'hbe1d1185), 
		.K5_C3_W0(32'hbd955177), .K5_C3_W1(32'hbdd5d39a), .K5_C3_W2(32'h3bb65b7e), .K5_C3_W3(32'hbdd48a75), .K5_C3_W4(32'hbd98c5fa), .K5_C3_W5(32'hbe12d82a), .K5_C3_W6(32'h3dc3e41b), .K5_C3_W7(32'hbe0a5dac), .K5_C3_W8(32'hbdad567f), 
		.K5_C4_W0(32'h3e3c0f83), .K5_C4_W1(32'hbdcdea92), .K5_C4_W2(32'h3e0f447c), .K5_C4_W3(32'h3d264e04), .K5_C4_W4(32'h3df884ad), .K5_C4_W5(32'h3de72ce7), .K5_C4_W6(32'hbdbf8dce), .K5_C4_W7(32'hbcdec684), .K5_C4_W8(32'hbdcef85d), 
		.K5_C5_W0(32'hbd6c166e), .K5_C5_W1(32'hbc87f2bd), .K5_C5_W2(32'hbd9bafc5), .K5_C5_W3(32'h3dff4527), .K5_C5_W4(32'h3e467462), .K5_C5_W5(32'hbdaac7f2), .K5_C5_W6(32'hbe25d7f4), .K5_C5_W7(32'hbbfdf75c), .K5_C5_W8(32'hbc466ae8), 
		.K5_C6_W0(32'hbd827093), .K5_C6_W1(32'hbc080025), .K5_C6_W2(32'h3de22d42), .K5_C6_W3(32'hbdd9340e), .K5_C6_W4(32'h3d4ccd32), .K5_C6_W5(32'h3b1a5820), .K5_C6_W6(32'hbd2944c0), .K5_C6_W7(32'hbc958072), .K5_C6_W8(32'hbe2e16bd), 
		.K5_C7_W0(32'hbe2a041f), .K5_C7_W1(32'h3de6a7e8), .K5_C7_W2(32'hbc3ae60d), .K5_C7_W3(32'hbdd4015e), .K5_C7_W4(32'h3d671a67), .K5_C7_W5(32'hbd85d9d8), .K5_C7_W6(32'h3c1b07e6), .K5_C7_W7(32'h3d6c282a), .K5_C7_W8(32'hbd96e66f), 
		.K5_BIAS (32'h3d0723d2),

		.K6_C0_W0(32'hbd58ad18), .K6_C0_W1(32'hbb9391fb), .K6_C0_W2(32'hbe1ae452), .K6_C0_W3(32'h3c6e5e5d), .K6_C0_W4(32'hba1e4b26), .K6_C0_W5(32'hbd9f8e23), .K6_C0_W6(32'hbce2bf48), .K6_C0_W7(32'h3e20b544), .K6_C0_W8(32'h3e10f556), 
		.K6_C1_W0(32'hbe1c4d3b), .K6_C1_W1(32'hbd26420d), .K6_C1_W2(32'h3cba98a6), .K6_C1_W3(32'h3d0e76bc), .K6_C1_W4(32'h3e2cb598), .K6_C1_W5(32'h3e092a57), .K6_C1_W6(32'hbe37ef88), .K6_C1_W7(32'hbd4c7f3b), .K6_C1_W8(32'h3e0fcc38), 
		.K6_C2_W0(32'hbcaf790e), .K6_C2_W1(32'h3d9745ef), .K6_C2_W2(32'h3e5b8807), .K6_C2_W3(32'hbd3795e5), .K6_C2_W4(32'h3dfa00a8), .K6_C2_W5(32'h3e33e2d5), .K6_C2_W6(32'hbdd87356), .K6_C2_W7(32'hbdf0d3a8), .K6_C2_W8(32'h3db0eb84), 
		.K6_C3_W0(32'h3dd4df79), .K6_C3_W1(32'hbe0966a6), .K6_C3_W2(32'h3d9e3ae0), .K6_C3_W3(32'hbe1e9d08), .K6_C3_W4(32'hbe16261b), .K6_C3_W5(32'h3e0110b4), .K6_C3_W6(32'hbcb1c787), .K6_C3_W7(32'h3d8fd2dc), .K6_C3_W8(32'h3de8389d), 
		.K6_C4_W0(32'h3de90ebf), .K6_C4_W1(32'h3dd3b86e), .K6_C4_W2(32'h3c9fe010), .K6_C4_W3(32'hbdf37cc1), .K6_C4_W4(32'hbdadbf30), .K6_C4_W5(32'hbdf1d908), .K6_C4_W6(32'hbd6a5415), .K6_C4_W7(32'h3d4ae819), .K6_C4_W8(32'hbe170255), 
		.K6_C5_W0(32'h3d0984c5), .K6_C5_W1(32'hbdc8b134), .K6_C5_W2(32'h3d06f584), .K6_C5_W3(32'h3d5980bd), .K6_C5_W4(32'h3d840fe9), .K6_C5_W5(32'h3df69448), .K6_C5_W6(32'h3da9cc39), .K6_C5_W7(32'h3da50cb0), .K6_C5_W8(32'hbd911512), 
		.K6_C6_W0(32'hbdc8cf5b), .K6_C6_W1(32'h3d85e0bf), .K6_C6_W2(32'hbb889de8), .K6_C6_W3(32'h3d18a557), .K6_C6_W4(32'hbb9301c9), .K6_C6_W5(32'hbc1565b5), .K6_C6_W6(32'h3d525984), .K6_C6_W7(32'h3cc9aed4), .K6_C6_W8(32'hbd12e78b), 
		.K6_C7_W0(32'hbd2671cc), .K6_C7_W1(32'h3af3f0a8), .K6_C7_W2(32'h3d80fe25), .K6_C7_W3(32'hbc8ab449), .K6_C7_W4(32'hbe1f80d4), .K6_C7_W5(32'hbdd26234), .K6_C7_W6(32'h3cec14ac), .K6_C7_W7(32'hbcd44810), .K6_C7_W8(32'hbd32521b), 
		.K6_BIAS (32'hbb0eeeee),

		.K7_C0_W0(32'hbdf81c76), .K7_C0_W1(32'h3de287eb), .K7_C0_W2(32'h3ce6bab9), .K7_C0_W3(32'hbdfc2d3f), .K7_C0_W4(32'hbd9bf7aa), .K7_C0_W5(32'hbdbff99e), .K7_C0_W6(32'h3b1c2e2d), .K7_C0_W7(32'hbd4e6808), .K7_C0_W8(32'hbccd62f0), 
		.K7_C1_W0(32'hbdb2ffe9), .K7_C1_W1(32'h3e1653d0), .K7_C1_W2(32'h3d851a72), .K7_C1_W3(32'h3dd92aa1), .K7_C1_W4(32'h3dcf62c0), .K7_C1_W5(32'hbdcc7de0), .K7_C1_W6(32'h3d659d14), .K7_C1_W7(32'h3e199414), .K7_C1_W8(32'hbd9f26e0), 
		.K7_C2_W0(32'hbe160723), .K7_C2_W1(32'h3e407372), .K7_C2_W2(32'hbdbdb8e9), .K7_C2_W3(32'hbc5d7b46), .K7_C2_W4(32'hbd4a86c5), .K7_C2_W5(32'h3e54fa2b), .K7_C2_W6(32'hbd99a51d), .K7_C2_W7(32'hbde6a2e5), .K7_C2_W8(32'h3e202577), 
		.K7_C3_W0(32'hbd7b8e8b), .K7_C3_W1(32'h3e024fa0), .K7_C3_W2(32'h3d8a1d0e), .K7_C3_W3(32'hbd81c84d), .K7_C3_W4(32'hbd84d3c4), .K7_C3_W5(32'h3d8d86d4), .K7_C3_W6(32'hbe00a4a8), .K7_C3_W7(32'hbd893cdc), .K7_C3_W8(32'h3e000676), 
		.K7_C4_W0(32'hbe12f2fa), .K7_C4_W1(32'hbd697bb1), .K7_C4_W2(32'h3e3df082), .K7_C4_W3(32'h3c3a6fc4), .K7_C4_W4(32'h3e2d488f), .K7_C4_W5(32'hbdd7840c), .K7_C4_W6(32'h3de4bf5d), .K7_C4_W7(32'h3e3ef070), .K7_C4_W8(32'hbdc8fec5), 
		.K7_C5_W0(32'hbd58ea49), .K7_C5_W1(32'hbdfca7e7), .K7_C5_W2(32'h3e337be2), .K7_C5_W3(32'hbe0840c9), .K7_C5_W4(32'hbe04c9c5), .K7_C5_W5(32'h3d2beead), .K7_C5_W6(32'h3d305400), .K7_C5_W7(32'h3cf9b88d), .K7_C5_W8(32'hbd57562e), 
		.K7_C6_W0(32'h3be41aae), .K7_C6_W1(32'hbdfa34c1), .K7_C6_W2(32'hbe249aed), .K7_C6_W3(32'h3e328679), .K7_C6_W4(32'h3b916702), .K7_C6_W5(32'h3dd52069), .K7_C6_W6(32'hbe313b1b), .K7_C6_W7(32'hbd9bbd21), .K7_C6_W8(32'hbd9b1aee), 
		.K7_C7_W0(32'hbe240bc2), .K7_C7_W1(32'hbdc028ea), .K7_C7_W2(32'hbd1dee37), .K7_C7_W3(32'h3d359fc0), .K7_C7_W4(32'h3dcf1f41), .K7_C7_W5(32'h3d9e6b77), .K7_C7_W6(32'h3e0f9a65), .K7_C7_W7(32'hbd0e250c), .K7_C7_W8(32'hbddf4eea), 
		.K7_BIAS (32'h3d5a813c),

		.K8_C0_W0(32'hbc8df81e), .K8_C0_W1(32'h3e276657), .K8_C0_W2(32'hbd231c97), .K8_C0_W3(32'hbe2ec898), .K8_C0_W4(32'h3e11ae1b), .K8_C0_W5(32'h3e013ebf), .K8_C0_W6(32'hbe2aed16), .K8_C0_W7(32'h3ca4ed72), .K8_C0_W8(32'h3d6f8dd8), 
		.K8_C1_W0(32'h3ddfdd75), .K8_C1_W1(32'hbe1a8584), .K8_C1_W2(32'hbd48d9fd), .K8_C1_W3(32'h3de76de5), .K8_C1_W4(32'hbd9bd974), .K8_C1_W5(32'h3e033e49), .K8_C1_W6(32'h3d98277e), .K8_C1_W7(32'hbb7ac556), .K8_C1_W8(32'h3cb33994), 
		.K8_C2_W0(32'hbd8b1ead), .K8_C2_W1(32'h3df0a41b), .K8_C2_W2(32'hbe50143f), .K8_C2_W3(32'hbe0599bb), .K8_C2_W4(32'h3db29513), .K8_C2_W5(32'h3dc25e77), .K8_C2_W6(32'hbe52510b), .K8_C2_W7(32'hbe45d4f2), .K8_C2_W8(32'h3d6568c3), 
		.K8_C3_W0(32'h3dca1753), .K8_C3_W1(32'h3dde53ad), .K8_C3_W2(32'h3ddea9f3), .K8_C3_W3(32'hbd183fff), .K8_C3_W4(32'h3d85b083), .K8_C3_W5(32'hbdaa02c1), .K8_C3_W6(32'hbd5404a6), .K8_C3_W7(32'h3c6b4ac6), .K8_C3_W8(32'h3e4099b7), 
		.K8_C4_W0(32'h3c9ed02b), .K8_C4_W1(32'h3d4b2e1e), .K8_C4_W2(32'hbd8f2211), .K8_C4_W3(32'hbe06aeca), .K8_C4_W4(32'hbd4e6823), .K8_C4_W5(32'h3e0ec14a), .K8_C4_W6(32'h3e1a1037), .K8_C4_W7(32'h3ddd1365), .K8_C4_W8(32'h3df48fa2), 
		.K8_C5_W0(32'h3d1db158), .K8_C5_W1(32'hbdd4e0ab), .K8_C5_W2(32'hbdbb6f6a), .K8_C5_W3(32'hbe2af1e4), .K8_C5_W4(32'hbdde72d5), .K8_C5_W5(32'hbd753f31), .K8_C5_W6(32'h3e08b468), .K8_C5_W7(32'h3e31213b), .K8_C5_W8(32'h3e1e6fe2), 
		.K8_C6_W0(32'hbddddf65), .K8_C6_W1(32'hbdd882df), .K8_C6_W2(32'h3e0fc638), .K8_C6_W3(32'h3e11d069), .K8_C6_W4(32'h3e0d1a01), .K8_C6_W5(32'hbdf070eb), .K8_C6_W6(32'h3d652722), .K8_C6_W7(32'hbe5ea9e4), .K8_C6_W8(32'hbd97aa20), 
		.K8_C7_W0(32'h3e3492a3), .K8_C7_W1(32'h3ddd2214), .K8_C7_W2(32'h3d8d9482), .K8_C7_W3(32'h3e5e4ed2), .K8_C7_W4(32'h3e02beb3), .K8_C7_W5(32'h3d2d8193), .K8_C7_W6(32'h3e3559c8), .K8_C7_W7(32'h3e034d14), .K8_C7_W8(32'h3e4b2fdd), 
		.K8_BIAS (32'hbcd436db),

		.K9_C0_W0(32'hbdac8109), .K9_C0_W1(32'hbe1df15a), .K9_C0_W2(32'hbe2591b5), .K9_C0_W3(32'hbae3f4f3), .K9_C0_W4(32'h3ce2202d), .K9_C0_W5(32'h3cec0668), .K9_C0_W6(32'h3dbdc7bb), .K9_C0_W7(32'h3d47f9c4), .K9_C0_W8(32'h3e29d86b), 
		.K9_C1_W0(32'h3e27535e), .K9_C1_W1(32'h3d9ca88b), .K9_C1_W2(32'hbe33af9f), .K9_C1_W3(32'hbdcbab21), .K9_C1_W4(32'hbd8d0765), .K9_C1_W5(32'hbe03c834), .K9_C1_W6(32'hbd696741), .K9_C1_W7(32'h3cff0b8e), .K9_C1_W8(32'hbe0df647), 
		.K9_C2_W0(32'hbcc78a5c), .K9_C2_W1(32'h3d03d5b8), .K9_C2_W2(32'h3e296425), .K9_C2_W3(32'h3da3d716), .K9_C2_W4(32'h3d922277), .K9_C2_W5(32'h3d5c9498), .K9_C2_W6(32'h3dd88748), .K9_C2_W7(32'h3e338afc), .K9_C2_W8(32'h3e45ca14), 
		.K9_C3_W0(32'h3d77e774), .K9_C3_W1(32'hbdb05569), .K9_C3_W2(32'h3e262892), .K9_C3_W3(32'hbdcd69ef), .K9_C3_W4(32'h3cf7275a), .K9_C3_W5(32'hbe24bda1), .K9_C3_W6(32'hbe1b4447), .K9_C3_W7(32'h3e18a0c8), .K9_C3_W8(32'h3d232e38), 
		.K9_C4_W0(32'hbd5e0fe8), .K9_C4_W1(32'hbdf4e7c7), .K9_C4_W2(32'hbcc7d809), .K9_C4_W3(32'hbc82914a), .K9_C4_W4(32'hba04b2c0), .K9_C4_W5(32'hbd7311d0), .K9_C4_W6(32'hba9359ab), .K9_C4_W7(32'h3d9b1f86), .K9_C4_W8(32'h3a9ecfc7), 
		.K9_C5_W0(32'h3d3f1f54), .K9_C5_W1(32'hbddc86f8), .K9_C5_W2(32'h3c543e2b), .K9_C5_W3(32'h3dad0002), .K9_C5_W4(32'hbd4cced9), .K9_C5_W5(32'h3dd6484c), .K9_C5_W6(32'h3e078411), .K9_C5_W7(32'hbe093400), .K9_C5_W8(32'h3e0e390a), 
		.K9_C6_W0(32'hbbdd2888), .K9_C6_W1(32'hbd510c33), .K9_C6_W2(32'hbdf3fcb9), .K9_C6_W3(32'h3d3641e5), .K9_C6_W4(32'h3e07edb4), .K9_C6_W5(32'h3dbeb3c8), .K9_C6_W6(32'hbd68a50e), .K9_C6_W7(32'h3e404d82), .K9_C6_W8(32'hbcd4224c), 
		.K9_C7_W0(32'hbe2714d2), .K9_C7_W1(32'hbe09bfa3), .K9_C7_W2(32'h3d7e71c7), .K9_C7_W3(32'hbdf5df71), .K9_C7_W4(32'h3d0f76dc), .K9_C7_W5(32'hbdde2aa1), .K9_C7_W6(32'hbdbdceba), .K9_C7_W7(32'h3ddc9fc1), .K9_C7_W8(32'hbd3503b4), 
		.K9_BIAS (32'h3cd2cbce),

		.K10_C0_W0(32'h3dc1c247), .K10_C0_W1(32'h3d5ce5b4), .K10_C0_W2(32'h3dbb0912), .K10_C0_W3(32'hbdbb9409), .K10_C0_W4(32'hbe1a5048), .K10_C0_W5(32'hbe08a0ee), .K10_C0_W6(32'hbe3630b6), .K10_C0_W7(32'hbd38214b), .K10_C0_W8(32'h3de5b5f5), 
		.K10_C1_W0(32'hbc646093), .K10_C1_W1(32'h3bba8afe), .K10_C1_W2(32'h3e4778fc), .K10_C1_W3(32'h3dccb5c5), .K10_C1_W4(32'h3d56fa63), .K10_C1_W5(32'hbcd7b8f2), .K10_C1_W6(32'hbd8e2a56), .K10_C1_W7(32'hbbb0fc3a), .K10_C1_W8(32'hbe112a6c), 
		.K10_C2_W0(32'hbc635e49), .K10_C2_W1(32'h3db43669), .K10_C2_W2(32'hbe361c2c), .K10_C2_W3(32'hbd99dac4), .K10_C2_W4(32'h3de8016b), .K10_C2_W5(32'h3e17723a), .K10_C2_W6(32'h3c8a7ffb), .K10_C2_W7(32'hbd730f81), .K10_C2_W8(32'hbd158bbb), 
		.K10_C3_W0(32'h3d140dcc), .K10_C3_W1(32'hbe2b01f9), .K10_C3_W2(32'hbbe9dc3e), .K10_C3_W3(32'hbe015542), .K10_C3_W4(32'hbd434a60), .K10_C3_W5(32'hbdbd9623), .K10_C3_W6(32'hbda11bae), .K10_C3_W7(32'h3e06e44b), .K10_C3_W8(32'hbdd95b34), 
		.K10_C4_W0(32'h3deb0f72), .K10_C4_W1(32'h3e0db731), .K10_C4_W2(32'hbce1fcee), .K10_C4_W3(32'hbd983224), .K10_C4_W4(32'hbd935e0d), .K10_C4_W5(32'h3e55a67c), .K10_C4_W6(32'hbdfe408b), .K10_C4_W7(32'h3e0703c1), .K10_C4_W8(32'h3d650cff), 
		.K10_C5_W0(32'h3df18351), .K10_C5_W1(32'h3de1079f), .K10_C5_W2(32'h3e35a239), .K10_C5_W3(32'h3d98392b), .K10_C5_W4(32'h3dd9adbd), .K10_C5_W5(32'h3ae22ced), .K10_C5_W6(32'hbe1ac940), .K10_C5_W7(32'hbdbd2989), .K10_C5_W8(32'hbdaadda4), 
		.K10_C6_W0(32'hbe05c9c5), .K10_C6_W1(32'h3d0388b0), .K10_C6_W2(32'hbd63aff3), .K10_C6_W3(32'hbd99b20e), .K10_C6_W4(32'h3d7e8b68), .K10_C6_W5(32'hbe07dba4), .K10_C6_W6(32'hbe53f59b), .K10_C6_W7(32'h3dba39e8), .K10_C6_W8(32'h3dc0c55f), 
		.K10_C7_W0(32'h3d97eaaa), .K10_C7_W1(32'h3d4e7363), .K10_C7_W2(32'hbd5fe99e), .K10_C7_W3(32'hbdccccb5), .K10_C7_W4(32'h3d468063), .K10_C7_W5(32'h3c2ea129), .K10_C7_W6(32'h3dbcb8cc), .K10_C7_W7(32'hbd8f3eab), .K10_C7_W8(32'hbe4c003c), 
		.K10_BIAS (32'h3cf2ccd2),

		.K11_C0_W0(32'hbd685ff4), .K11_C0_W1(32'h3d93b49b), .K11_C0_W2(32'h3e2b957a), .K11_C0_W3(32'h3d182bbb), .K11_C0_W4(32'h3c513b12), .K11_C0_W5(32'hbdafb57a), .K11_C0_W6(32'hbcff9e66), .K11_C0_W7(32'h3c88a1c5), .K11_C0_W8(32'hbce2e039), 
		.K11_C1_W0(32'hbd003b2a), .K11_C1_W1(32'hbe18d07c), .K11_C1_W2(32'hbc9f8075), .K11_C1_W3(32'h3c2c7cbc), .K11_C1_W4(32'hbce1e185), .K11_C1_W5(32'hbdb6776b), .K11_C1_W6(32'h3d6a132f), .K11_C1_W7(32'h3e191809), .K11_C1_W8(32'h3e1f0eb3), 
		.K11_C2_W0(32'hbdedf09c), .K11_C2_W1(32'h3defc5e0), .K11_C2_W2(32'hbc1fda1b), .K11_C2_W3(32'hbe15b1f9), .K11_C2_W4(32'hbc27cd63), .K11_C2_W5(32'h3dd91534), .K11_C2_W6(32'hbd1e34b1), .K11_C2_W7(32'h3d0fd199), .K11_C2_W8(32'hb9f1e1c8), 
		.K11_C3_W0(32'h3e320b47), .K11_C3_W1(32'h3d98decc), .K11_C3_W2(32'hbd081839), .K11_C3_W3(32'h3d1c1ecc), .K11_C3_W4(32'h3dbf7409), .K11_C3_W5(32'hbe1349e2), .K11_C3_W6(32'hbc5119b1), .K11_C3_W7(32'hbdc9cc8a), .K11_C3_W8(32'hbd9c603d), 
		.K11_C4_W0(32'hbd828791), .K11_C4_W1(32'hbd94ab28), .K11_C4_W2(32'hbe2058d3), .K11_C4_W3(32'h3e2339d4), .K11_C4_W4(32'h3da2c135), .K11_C4_W5(32'hbe0d1210), .K11_C4_W6(32'hbdd7ae21), .K11_C4_W7(32'h3da1c651), .K11_C4_W8(32'hbda651ab), 
		.K11_C5_W0(32'h3d85a49e), .K11_C5_W1(32'hbdd0ff3e), .K11_C5_W2(32'hbd727f8d), .K11_C5_W3(32'hbe15d260), .K11_C5_W4(32'h3e05727f), .K11_C5_W5(32'h3e0f62dd), .K11_C5_W6(32'hbd740511), .K11_C5_W7(32'hbe070936), .K11_C5_W8(32'h3c9d0f36), 
		.K11_C6_W0(32'h3e0f06db), .K11_C6_W1(32'hbc4a15ae), .K11_C6_W2(32'hbde9ed83), .K11_C6_W3(32'hbd8e7430), .K11_C6_W4(32'hbd91721a), .K11_C6_W5(32'h3e08c43e), .K11_C6_W6(32'h3e12ba0d), .K11_C6_W7(32'hbe1978f7), .K11_C6_W8(32'h3c2c4cac), 
		.K11_C7_W0(32'h3d33bec6), .K11_C7_W1(32'h3dbe0e19), .K11_C7_W2(32'h3da84853), .K11_C7_W3(32'h3dd8af3e), .K11_C7_W4(32'h3e282cc2), .K11_C7_W5(32'hbcaa053a), .K11_C7_W6(32'hbd478e03), .K11_C7_W7(32'hbde0bb6e), .K11_C7_W8(32'h3df39801), 
		.K11_BIAS (32'hbc93f8d3),

		.K12_C0_W0(32'h3d1cf06f), .K12_C0_W1(32'hbd8829ea), .K12_C0_W2(32'hbc8f0065), .K12_C0_W3(32'hbd86ba70), .K12_C0_W4(32'h3d6187d8), .K12_C0_W5(32'hba34a764), .K12_C0_W6(32'h3dd24465), .K12_C0_W7(32'h3dc132f7), .K12_C0_W8(32'hbb37af59), 
		.K12_C1_W0(32'hbc400d0d), .K12_C1_W1(32'hbd1c4d66), .K12_C1_W2(32'hbd12a334), .K12_C1_W3(32'h3dacb923), .K12_C1_W4(32'h3c2a6f57), .K12_C1_W5(32'h3dc49d8a), .K12_C1_W6(32'h3e0525e8), .K12_C1_W7(32'h3df79a6a), .K12_C1_W8(32'hbdb7fd13), 
		.K12_C2_W0(32'h3e775491), .K12_C2_W1(32'h3d8707ea), .K12_C2_W2(32'hbdb55214), .K12_C2_W3(32'h3c8333c7), .K12_C2_W4(32'h39d31e96), .K12_C2_W5(32'hbe25a6ed), .K12_C2_W6(32'hbc0b535b), .K12_C2_W7(32'hbde174c2), .K12_C2_W8(32'h3dc4d6d3), 
		.K12_C3_W0(32'h3e27887c), .K12_C3_W1(32'h3e394561), .K12_C3_W2(32'hbd461ff2), .K12_C3_W3(32'hbd9d85fc), .K12_C3_W4(32'h3e1febc9), .K12_C3_W5(32'hbd688658), .K12_C3_W6(32'h3d847b6e), .K12_C3_W7(32'h3d0d89db), .K12_C3_W8(32'h3db344a1), 
		.K12_C4_W0(32'hbe07611c), .K12_C4_W1(32'h3df599ce), .K12_C4_W2(32'hbd88850f), .K12_C4_W3(32'h3db67f83), .K12_C4_W4(32'hbe353bb8), .K12_C4_W5(32'h3c1002be), .K12_C4_W6(32'hbd408acc), .K12_C4_W7(32'h3c5d6de3), .K12_C4_W8(32'hbce4907d), 
		.K12_C5_W0(32'h3d8abb41), .K12_C5_W1(32'hbe0f0143), .K12_C5_W2(32'hbd67eaf9), .K12_C5_W3(32'h3daf59c9), .K12_C5_W4(32'h3de1b855), .K12_C5_W5(32'hbc652f41), .K12_C5_W6(32'h3dd4c7ee), .K12_C5_W7(32'h3d858d22), .K12_C5_W8(32'hbcd769f0), 
		.K12_C6_W0(32'hbcf8918e), .K12_C6_W1(32'h3be71e71), .K12_C6_W2(32'h3e3cc499), .K12_C6_W3(32'h3d4ca24d), .K12_C6_W4(32'h3e1ba8c9), .K12_C6_W5(32'h3e387a9e), .K12_C6_W6(32'hbe44e7f9), .K12_C6_W7(32'hbe4fd78e), .K12_C6_W8(32'hbe318969), 
		.K12_C7_W0(32'hbe0c8f86), .K12_C7_W1(32'hbd10c746), .K12_C7_W2(32'h3da4a368), .K12_C7_W3(32'h3d07ccad), .K12_C7_W4(32'h3c556923), .K12_C7_W5(32'h3cf77eaf), .K12_C7_W6(32'h3c78c91f), .K12_C7_W7(32'h3dd7b450), .K12_C7_W8(32'hbe09e6f7), 
		.K12_BIAS (32'hbcf530be),

		.K13_C0_W0(32'h3e04a90e), .K13_C0_W1(32'h3cb04d94), .K13_C0_W2(32'hbe0980fb), .K13_C0_W3(32'h3e07e8ba), .K13_C0_W4(32'h3e282673), .K13_C0_W5(32'h3e008992), .K13_C0_W6(32'hbdb93be4), .K13_C0_W7(32'h3d906541), .K13_C0_W8(32'h3da192ad), 
		.K13_C1_W0(32'hbdf500a3), .K13_C1_W1(32'hbd9044cf), .K13_C1_W2(32'hbd446db1), .K13_C1_W3(32'hbdce905a), .K13_C1_W4(32'h3d4111a8), .K13_C1_W5(32'h3d643a12), .K13_C1_W6(32'hbdf93d23), .K13_C1_W7(32'h3d4e9d29), .K13_C1_W8(32'hbbe26aa3), 
		.K13_C2_W0(32'hbd54477a), .K13_C2_W1(32'hbe2c7a44), .K13_C2_W2(32'h3d6967cf), .K13_C2_W3(32'hbdad6e88), .K13_C2_W4(32'hbd25697a), .K13_C2_W5(32'h3db634bd), .K13_C2_W6(32'h3d0f3d31), .K13_C2_W7(32'hbe2019ad), .K13_C2_W8(32'hbd8b5af2), 
		.K13_C3_W0(32'h3e06fed5), .K13_C3_W1(32'h3e032ca6), .K13_C3_W2(32'hbd4de381), .K13_C3_W3(32'hbd86e865), .K13_C3_W4(32'h3d23339f), .K13_C3_W5(32'hbdcef961), .K13_C3_W6(32'hbd67e807), .K13_C3_W7(32'h3d2f375e), .K13_C3_W8(32'h3e28c31b), 
		.K13_C4_W0(32'h3d59c91b), .K13_C4_W1(32'hbe0b17fd), .K13_C4_W2(32'h3b10c1fa), .K13_C4_W3(32'hbdee6c7c), .K13_C4_W4(32'hbd8aed31), .K13_C4_W5(32'hbc668c4b), .K13_C4_W6(32'hbdbc7068), .K13_C4_W7(32'hbe094552), .K13_C4_W8(32'h3e2bc0b4), 
		.K13_C5_W0(32'h3e1b650e), .K13_C5_W1(32'h3ddbac99), .K13_C5_W2(32'h3d8b9794), .K13_C5_W3(32'hbd83eeb7), .K13_C5_W4(32'h3e2fa336), .K13_C5_W5(32'hbd641adc), .K13_C5_W6(32'hbd351018), .K13_C5_W7(32'h3e20b6f4), .K13_C5_W8(32'h3e038fdf), 
		.K13_C6_W0(32'hbe148228), .K13_C6_W1(32'hbdc80a85), .K13_C6_W2(32'hbd8f4fd4), .K13_C6_W3(32'h3e3702dd), .K13_C6_W4(32'h3dd44011), .K13_C6_W5(32'hbcc793f4), .K13_C6_W6(32'h3dfd9a34), .K13_C6_W7(32'h3d2a53f6), .K13_C6_W8(32'hbd44a8ff), 
		.K13_C7_W0(32'hbc848907), .K13_C7_W1(32'hba7ec877), .K13_C7_W2(32'h3d809df0), .K13_C7_W3(32'h3e1f3e17), .K13_C7_W4(32'hbd9b2b87), .K13_C7_W5(32'hbd938e1e), .K13_C7_W6(32'hbd26d658), .K13_C7_W7(32'hbdee2819), .K13_C7_W8(32'h3c518970), 
		.K13_BIAS (32'hbceec530),

		.K14_C0_W0(32'hbdf1a440), .K14_C0_W1(32'h3dacd125), .K14_C0_W2(32'h3e1c4c7a), .K14_C0_W3(32'h3e18c184), .K14_C0_W4(32'hbe0c77d0), .K14_C0_W5(32'hbccffbfe), .K14_C0_W6(32'h3e3f497c), .K14_C0_W7(32'hbe1a0f3a), .K14_C0_W8(32'hbddb6518), 
		.K14_C1_W0(32'hbdca28d3), .K14_C1_W1(32'h3d9becdb), .K14_C1_W2(32'h3dfae6f9), .K14_C1_W3(32'hbc95fb69), .K14_C1_W4(32'h3c486c05), .K14_C1_W5(32'h3d44e84f), .K14_C1_W6(32'hbe26149b), .K14_C1_W7(32'h3c85d0bd), .K14_C1_W8(32'h3dcb2f32), 
		.K14_C2_W0(32'hbdc5aa96), .K14_C2_W1(32'hbe07352e), .K14_C2_W2(32'hbd37c5ae), .K14_C2_W3(32'h3d5c29ca), .K14_C2_W4(32'hbe0e0bb8), .K14_C2_W5(32'hbde89807), .K14_C2_W6(32'hbcc7cd1f), .K14_C2_W7(32'hbd2035bd), .K14_C2_W8(32'h3d281798), 
		.K14_C3_W0(32'hbd49f8d0), .K14_C3_W1(32'hbd34af31), .K14_C3_W2(32'h3e0af9ff), .K14_C3_W3(32'hbdc81ab7), .K14_C3_W4(32'hbdbb9277), .K14_C3_W5(32'hbd51d4e8), .K14_C3_W6(32'h3da57fdd), .K14_C3_W7(32'hbceafe0c), .K14_C3_W8(32'hbda2e9d3), 
		.K14_C4_W0(32'hbe1fcafc), .K14_C4_W1(32'h3d9329fe), .K14_C4_W2(32'hbd6f8a98), .K14_C4_W3(32'hbe2e0a75), .K14_C4_W4(32'hbe09016f), .K14_C4_W5(32'hbc44a5c2), .K14_C4_W6(32'h3a41c5ac), .K14_C4_W7(32'hbcbdf369), .K14_C4_W8(32'h3e307ef1), 
		.K14_C5_W0(32'h3d3deb57), .K14_C5_W1(32'hbdccdce5), .K14_C5_W2(32'h3dfb047e), .K14_C5_W3(32'hbe07ae39), .K14_C5_W4(32'h3d8f0233), .K14_C5_W5(32'hbdf8d611), .K14_C5_W6(32'hbe325a9f), .K14_C5_W7(32'h3cafda71), .K14_C5_W8(32'hbe2094c0), 
		.K14_C6_W0(32'hbe1a10be), .K14_C6_W1(32'h3ca7eb74), .K14_C6_W2(32'hbe2b2a79), .K14_C6_W3(32'h3d50bd02), .K14_C6_W4(32'hbcc8976f), .K14_C6_W5(32'h3dee2e29), .K14_C6_W6(32'hbd0f504d), .K14_C6_W7(32'hbd951e5a), .K14_C6_W8(32'hbd0c3336), 
		.K14_C7_W0(32'hbe22821b), .K14_C7_W1(32'h3d998dff), .K14_C7_W2(32'h3d846192), .K14_C7_W3(32'h3d2e28ab), .K14_C7_W4(32'h3e38bf17), .K14_C7_W5(32'h3e3e0cc3), .K14_C7_W6(32'h3d7fc125), .K14_C7_W7(32'hbcb2d319), .K14_C7_W8(32'h3e00eea7), 
		.K14_BIAS (32'hbb80d1f9),

		.K15_C0_W0(32'h3dc06f78), .K15_C0_W1(32'h3dcdf944), .K15_C0_W2(32'h3daf3151), .K15_C0_W3(32'h3de11fa7), .K15_C0_W4(32'h3dd20359), .K15_C0_W5(32'hbd212509), .K15_C0_W6(32'hbdf60245), .K15_C0_W7(32'h3df53491), .K15_C0_W8(32'hbdd51628), 
		.K15_C1_W0(32'hbd14fa24), .K15_C1_W1(32'hbd93b814), .K15_C1_W2(32'hbdc5317e), .K15_C1_W3(32'h3e257438), .K15_C1_W4(32'hbd003158), .K15_C1_W5(32'hbcda0b86), .K15_C1_W6(32'h3c72e4dd), .K15_C1_W7(32'h3dabfc98), .K15_C1_W8(32'h3dfe3bdb), 
		.K15_C2_W0(32'h3d298831), .K15_C2_W1(32'hbd67c0e2), .K15_C2_W2(32'hbb1d47be), .K15_C2_W3(32'h3dc62134), .K15_C2_W4(32'hbdf1d0d5), .K15_C2_W5(32'hbdf56b9f), .K15_C2_W6(32'h3d09f5ea), .K15_C2_W7(32'hbe39b131), .K15_C2_W8(32'hbe201dbc), 
		.K15_C3_W0(32'h3e07adb3), .K15_C3_W1(32'hbda5ba6f), .K15_C3_W2(32'hbb56baad), .K15_C3_W3(32'hbd0009d2), .K15_C3_W4(32'h3e1abdd9), .K15_C3_W5(32'h3e5e8210), .K15_C3_W6(32'h3d5d7a2c), .K15_C3_W7(32'hbe0f9d17), .K15_C3_W8(32'hbde10488), 
		.K15_C4_W0(32'hbe1fbc7c), .K15_C4_W1(32'h3e20f11b), .K15_C4_W2(32'hbdc2f4ef), .K15_C4_W3(32'h3d1759a6), .K15_C4_W4(32'h3e2dfc7d), .K15_C4_W5(32'hbc608175), .K15_C4_W6(32'hbd46ad0f), .K15_C4_W7(32'h3d79c35b), .K15_C4_W8(32'hbdedd9e4), 
		.K15_C5_W0(32'h3e187ed1), .K15_C5_W1(32'hbde28e1b), .K15_C5_W2(32'hbd91a009), .K15_C5_W3(32'hbd9a462e), .K15_C5_W4(32'h3e052989), .K15_C5_W5(32'hbdc39c38), .K15_C5_W6(32'h3d9ab74a), .K15_C5_W7(32'h3e3cadaa), .K15_C5_W8(32'h3d84825d), 
		.K15_C6_W0(32'hbd97cb24), .K15_C6_W1(32'hbe0756f4), .K15_C6_W2(32'hbd9e2bde), .K15_C6_W3(32'hbda3bc12), .K15_C6_W4(32'hbe0d65ee), .K15_C6_W5(32'hbda346b2), .K15_C6_W6(32'hbc97eb80), .K15_C6_W7(32'hbcb785ba), .K15_C6_W8(32'hbb98da6a), 
		.K15_C7_W0(32'h3c827f28), .K15_C7_W1(32'hbac4a192), .K15_C7_W2(32'h3db778cd), .K15_C7_W3(32'hbd2313c6), .K15_C7_W4(32'h3d86816c), .K15_C7_W5(32'h3e20a0a3), .K15_C7_W6(32'hbe1d8f95), .K15_C7_W7(32'h3e3a3eaf), .K15_C7_W8(32'hbc60d034), 
		.K15_BIAS (32'h3c3d7ea9)
		)
		block4_conv1(
		.clk(clk),
		.resetn(resetn),
		.data_valid_in(valid_in),
		.data_in_0(data_in_0),
		.data_in_1(data_in_1),
		.data_in_2(data_in_2),
		.data_in_3(data_in_3),
		.data_in_4(data_in_4),
		.data_in_5(data_in_5),
		.data_in_6(data_in_6),
		.data_in_7(data_in_7),
		.data_out_conv_0(conv_out_4_1[0]),
		.data_out_conv_1(conv_out_4_1[1]),
		.data_out_conv_2(conv_out_4_1[2]),
		.data_out_conv_3(conv_out_4_1[3]),
		.data_out_conv_4(conv_out_4_1[4]),
		.data_out_conv_5(conv_out_4_1[5]),
		.data_out_conv_6(conv_out_4_1[6]),
		.data_out_conv_7(conv_out_4_1[7]),
		.data_out_conv_8(conv_out_4_1[8]),
		.data_out_conv_9(conv_out_4_1[9]),
		.data_out_conv_10(conv_out_4_1[10]),
		.data_out_conv_11(conv_out_4_1[11]),
		.data_out_conv_12(conv_out_4_1[12]),
		.data_out_conv_13(conv_out_4_1[13]),
		.data_out_conv_14(conv_out_4_1[14]),
		.data_out_conv_15(conv_out_4_1[15]),
		.valid_out_pixel(conv_valid_out_4_1),
		.done(done_conv_4_1)
		);   





	conv3d_16_kernel_16_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(WIDTH),.IMG_HEIGHT(HEIGHT),
		.K0_C0_W0(32'h3db42524), .K0_C0_W1(32'hbe137928), .K0_C0_W2(32'h3cb68062), .K0_C0_W3(32'hbe2091d5), .K0_C0_W4(32'hbd927ef5), .K0_C0_W5(32'h3de56c8a), .K0_C0_W6(32'h3c841ece), .K0_C0_W7(32'h3c98ae5b), .K0_C0_W8(32'hbd67f492), 
		.K0_C1_W0(32'hbd975271), .K0_C1_W1(32'hbd13fb91), .K0_C1_W2(32'h3ddab69a), .K0_C1_W3(32'h3df50350), .K0_C1_W4(32'hbddf3c8e), .K0_C1_W5(32'h3db9e3d5), .K0_C1_W6(32'hbb67b877), .K0_C1_W7(32'hbd9bf183), .K0_C1_W8(32'h3e15f132), 
		.K0_C2_W0(32'hbe0d012d), .K0_C2_W1(32'hbd0bf445), .K0_C2_W2(32'hbde408db), .K0_C2_W3(32'h3c87e623), .K0_C2_W4(32'hbd32f11f), .K0_C2_W5(32'h3c6938c6), .K0_C2_W6(32'hbdf4798f), .K0_C2_W7(32'h3d265b34), .K0_C2_W8(32'h3d64ecf9), 
		.K0_C3_W0(32'hbccfa8d3), .K0_C3_W1(32'h3b1f7ea5), .K0_C3_W2(32'hbd6d915d), .K0_C3_W3(32'hbdc26561), .K0_C3_W4(32'hbd8721c8), .K0_C3_W5(32'h3dbcf23b), .K0_C3_W6(32'h3da9e268), .K0_C3_W7(32'hbdbffdbc), .K0_C3_W8(32'hbe096088), 
		.K0_C4_W0(32'h3d71083c), .K0_C4_W1(32'hbdd08959), .K0_C4_W2(32'hbc439d7c), .K0_C4_W3(32'hbe11beb8), .K0_C4_W4(32'h3d9abf7f), .K0_C4_W5(32'h3dcf164b), .K0_C4_W6(32'h3c162d34), .K0_C4_W7(32'h3e0c9a16), .K0_C4_W8(32'hbde897d0), 
		.K0_C5_W0(32'h3d973355), .K0_C5_W1(32'hbddd6cb8), .K0_C5_W2(32'h3d0090ba), .K0_C5_W3(32'h3e191ec4), .K0_C5_W4(32'h3e1964d9), .K0_C5_W5(32'hbd4c19ad), .K0_C5_W6(32'h3caa4183), .K0_C5_W7(32'hbd7de357), .K0_C5_W8(32'hbdd3d730), 
		.K0_C6_W0(32'hbac9fcc7), .K0_C6_W1(32'hbd7d441d), .K0_C6_W2(32'h3b2654bc), .K0_C6_W3(32'hbd0232fb), .K0_C6_W4(32'hbd32b25e), .K0_C6_W5(32'h3de6e41d), .K0_C6_W6(32'hbdb5f28c), .K0_C6_W7(32'hbcc1fc7c), .K0_C6_W8(32'h3d997f5f), 
		.K0_C7_W0(32'h3cdaace6), .K0_C7_W1(32'h3dac4377), .K0_C7_W2(32'h3d45ee25), .K0_C7_W3(32'hbd4240ad), .K0_C7_W4(32'h3cf9ee14), .K0_C7_W5(32'hbe0527c9), .K0_C7_W6(32'h3d366eb4), .K0_C7_W7(32'h3dba649f), .K0_C7_W8(32'hbdee128b), 
		.K0_C8_W0(32'hbbd561be), .K0_C8_W1(32'hbdd64a39), .K0_C8_W2(32'h3e014958), .K0_C8_W3(32'h3cb227e0), .K0_C8_W4(32'hbded85f9), .K0_C8_W5(32'h3dbe3ca6), .K0_C8_W6(32'hbdfae2d6), .K0_C8_W7(32'h3d1f63b0), .K0_C8_W8(32'h3d84d082), 
		.K0_C9_W0(32'hbdc73eab), .K0_C9_W1(32'h3db139d3), .K0_C9_W2(32'h3cee2b4a), .K0_C9_W3(32'hbdfae943), .K0_C9_W4(32'hbdafd917), .K0_C9_W5(32'hbdb7790f), .K0_C9_W6(32'hbc9da99c), .K0_C9_W7(32'hbb8c7306), .K0_C9_W8(32'hbde26914), 
		.K0_C10_W0(32'hbddf25af), .K0_C10_W1(32'hbd067c76), .K0_C10_W2(32'hbdbc901d), .K0_C10_W3(32'hb9e637cd), .K0_C10_W4(32'h3c854457), .K0_C10_W5(32'h3d43eff1), .K0_C10_W6(32'h3d46838c), .K0_C10_W7(32'h3d96de4f), .K0_C10_W8(32'h3d4733a0), 
		.K0_C11_W0(32'h3e0fd04b), .K0_C11_W1(32'h3daf4b78), .K0_C11_W2(32'hbca87aee), .K0_C11_W3(32'hbaa5aa79), .K0_C11_W4(32'hbc5173e7), .K0_C11_W5(32'h3da90185), .K0_C11_W6(32'h3da7edee), .K0_C11_W7(32'hbcfafb0a), .K0_C11_W8(32'hbd4ebb57), 
		.K0_C12_W0(32'h3e1bd117), .K0_C12_W1(32'h3dcadb0c), .K0_C12_W2(32'h3de994e4), .K0_C12_W3(32'hbd8c3458), .K0_C12_W4(32'h3d5fe752), .K0_C12_W5(32'h3e131da8), .K0_C12_W6(32'hbcf605e1), .K0_C12_W7(32'h3ba4e8eb), .K0_C12_W8(32'hbe0f6a10), 
		.K0_C13_W0(32'hbe117fe4), .K0_C13_W1(32'hbd231651), .K0_C13_W2(32'h3d671e6b), .K0_C13_W3(32'hbc51d5f0), .K0_C13_W4(32'hbe0ad761), .K0_C13_W5(32'hbd1619d6), .K0_C13_W6(32'hbe199ec5), .K0_C13_W7(32'h3ca17876), .K0_C13_W8(32'hbdc81da9), 
		.K0_C14_W0(32'hbddaaeb4), .K0_C14_W1(32'hbcf83d15), .K0_C14_W2(32'hbc662459), .K0_C14_W3(32'hbc649c3f), .K0_C14_W4(32'hbde5e8bb), .K0_C14_W5(32'hbc94500b), .K0_C14_W6(32'h3dc23112), .K0_C14_W7(32'hbc5aa234), .K0_C14_W8(32'h3c15340f), 
		.K0_C15_W0(32'hbc67b69a), .K0_C15_W1(32'h3d8cbdfb), .K0_C15_W2(32'hbdc24bfb), .K0_C15_W3(32'h3dda5ab6), .K0_C15_W4(32'hbaedb720), .K0_C15_W5(32'hbda2b0e4), .K0_C15_W6(32'h3cee3fc8), .K0_C15_W7(32'hbc65974b), .K0_C15_W8(32'h3d86e83b), 
		.K0_BIAS (32'h3ca0475d),

		.K1_C0_W0(32'h3e03f1f2), .K1_C0_W1(32'hbe0824d3), .K1_C0_W2(32'hbe3058d6), .K1_C0_W3(32'hbde21627), .K1_C0_W4(32'hbd17a0e3), .K1_C0_W5(32'hbda5ca14), .K1_C0_W6(32'hbe0000c1), .K1_C0_W7(32'hbacfe0cc), .K1_C0_W8(32'h3b8efb29), 
		.K1_C1_W0(32'h3c25141b), .K1_C1_W1(32'h3d691403), .K1_C1_W2(32'h3d0d614f), .K1_C1_W3(32'h3e04bf56), .K1_C1_W4(32'hbd813449), .K1_C1_W5(32'h3d31e387), .K1_C1_W6(32'hbddaccd7), .K1_C1_W7(32'hbde5a95f), .K1_C1_W8(32'h3d4974a4), 
		.K1_C2_W0(32'h3e06a862), .K1_C2_W1(32'h3bf5b250), .K1_C2_W2(32'hbdfec480), .K1_C2_W3(32'h3de923c5), .K1_C2_W4(32'h3bc7eba0), .K1_C2_W5(32'hbddeb2f2), .K1_C2_W6(32'hbd825740), .K1_C2_W7(32'hbdefcba2), .K1_C2_W8(32'h3d3cd8fc), 
		.K1_C3_W0(32'hbbd1824c), .K1_C3_W1(32'h3d114910), .K1_C3_W2(32'h3df575b2), .K1_C3_W3(32'h3de42c95), .K1_C3_W4(32'h3d899d09), .K1_C3_W5(32'h3e04972c), .K1_C3_W6(32'hbdf92033), .K1_C3_W7(32'hbdeba4dd), .K1_C3_W8(32'h3b7002d5), 
		.K1_C4_W0(32'h3c1c45f0), .K1_C4_W1(32'hbbbc8358), .K1_C4_W2(32'h3db6669f), .K1_C4_W3(32'hbdf95d6b), .K1_C4_W4(32'h3ca529af), .K1_C4_W5(32'hbe04bb03), .K1_C4_W6(32'hbd74e315), .K1_C4_W7(32'h3cad589d), .K1_C4_W8(32'hbde476f4), 
		.K1_C5_W0(32'h3df62d65), .K1_C5_W1(32'h3db79f9c), .K1_C5_W2(32'h3cd7ec34), .K1_C5_W3(32'h3d08442a), .K1_C5_W4(32'h3daaa97d), .K1_C5_W5(32'h3d366e45), .K1_C5_W6(32'h3962b188), .K1_C5_W7(32'hbd22b433), .K1_C5_W8(32'h3da5bba0), 
		.K1_C6_W0(32'h3cdd2c27), .K1_C6_W1(32'hbd5306f2), .K1_C6_W2(32'hbd9fbac9), .K1_C6_W3(32'h3d1662fc), .K1_C6_W4(32'h3d4ed406), .K1_C6_W5(32'h3cfc6d09), .K1_C6_W6(32'hbd92b152), .K1_C6_W7(32'hbdada4c9), .K1_C6_W8(32'hbd4cf682), 
		.K1_C7_W0(32'h3c2ab086), .K1_C7_W1(32'h3e18e091), .K1_C7_W2(32'h3dead7ad), .K1_C7_W3(32'h3cd6f99d), .K1_C7_W4(32'hbcc4a8ec), .K1_C7_W5(32'h3d9f3e44), .K1_C7_W6(32'hbe08b5fc), .K1_C7_W7(32'h3dfff981), .K1_C7_W8(32'hbdf6f37f), 
		.K1_C8_W0(32'h3d562bbb), .K1_C8_W1(32'h3c2ec47d), .K1_C8_W2(32'h3e08370d), .K1_C8_W3(32'hbcaabc8d), .K1_C8_W4(32'h3d57d799), .K1_C8_W5(32'h3ce0768e), .K1_C8_W6(32'hbdcb81fe), .K1_C8_W7(32'hbdc9c339), .K1_C8_W8(32'h3d85ccbf), 
		.K1_C9_W0(32'hbdd15ac3), .K1_C9_W1(32'h3d924a19), .K1_C9_W2(32'hbd234360), .K1_C9_W3(32'h3e1ec250), .K1_C9_W4(32'h3e01f0a4), .K1_C9_W5(32'hbe0acc3e), .K1_C9_W6(32'hbdea7b95), .K1_C9_W7(32'hbcf0cf5b), .K1_C9_W8(32'hbd87747e), 
		.K1_C10_W0(32'h3ce64554), .K1_C10_W1(32'h3dfcbf6c), .K1_C10_W2(32'h3b83fa8d), .K1_C10_W3(32'hbde5e324), .K1_C10_W4(32'h3cedb27a), .K1_C10_W5(32'h3c7b5e10), .K1_C10_W6(32'h3ce83a75), .K1_C10_W7(32'hbda84f1a), .K1_C10_W8(32'h3e047c76), 
		.K1_C11_W0(32'hbded9dcb), .K1_C11_W1(32'hbd25c49c), .K1_C11_W2(32'hbde935d9), .K1_C11_W3(32'h3d1df2f5), .K1_C11_W4(32'h3e1d1fce), .K1_C11_W5(32'h3c6929b0), .K1_C11_W6(32'hbe1a26be), .K1_C11_W7(32'hbd6239d6), .K1_C11_W8(32'h3bfb5871), 
		.K1_C12_W0(32'h3db10a89), .K1_C12_W1(32'hbddef42f), .K1_C12_W2(32'hbdd11aa3), .K1_C12_W3(32'h3d87e9ee), .K1_C12_W4(32'hbc85fea5), .K1_C12_W5(32'h3ceffd2a), .K1_C12_W6(32'hbc0f98d2), .K1_C12_W7(32'hbde64718), .K1_C12_W8(32'h3d178f08), 
		.K1_C13_W0(32'h3dfa73fa), .K1_C13_W1(32'h3dc4abbd), .K1_C13_W2(32'h3d79bf8c), .K1_C13_W3(32'hbd589d97), .K1_C13_W4(32'hbd71cf27), .K1_C13_W5(32'hbd5655fc), .K1_C13_W6(32'hbcf00dcf), .K1_C13_W7(32'hbdfab526), .K1_C13_W8(32'h3d7ee223), 
		.K1_C14_W0(32'hbd561503), .K1_C14_W1(32'hbd97c9ab), .K1_C14_W2(32'hbcd83b50), .K1_C14_W3(32'h3dc9f8ad), .K1_C14_W4(32'h3cb1adcc), .K1_C14_W5(32'hbd85c13c), .K1_C14_W6(32'hbdcad0cb), .K1_C14_W7(32'hbdd3ffd8), .K1_C14_W8(32'h3d5730d2), 
		.K1_C15_W0(32'hbdd9c548), .K1_C15_W1(32'hbd4623f1), .K1_C15_W2(32'hbe0d6ff5), .K1_C15_W3(32'hbce272e8), .K1_C15_W4(32'h3c21b727), .K1_C15_W5(32'h3d33319c), .K1_C15_W6(32'hbdb770bf), .K1_C15_W7(32'hbd1d9895), .K1_C15_W8(32'hbba7dad0), 
		.K1_BIAS (32'hbc007778),

		.K2_C0_W0(32'h3e0d6a66), .K2_C0_W1(32'h3d5db55f), .K2_C0_W2(32'h3d8d348e), .K2_C0_W3(32'h3d03c93c), .K2_C0_W4(32'hbdb228b9), .K2_C0_W5(32'h3d699555), .K2_C0_W6(32'h3cb4b7fd), .K2_C0_W7(32'hbccb8d83), .K2_C0_W8(32'h3e027439), 
		.K2_C1_W0(32'hbc219ecc), .K2_C1_W1(32'h3cf829ab), .K2_C1_W2(32'h3dce43b1), .K2_C1_W3(32'hbddac4ae), .K2_C1_W4(32'hbbc5a772), .K2_C1_W5(32'h3de858b7), .K2_C1_W6(32'hbaf88183), .K2_C1_W7(32'h3d78da5a), .K2_C1_W8(32'h3e08543d), 
		.K2_C2_W0(32'hbd0ccd3b), .K2_C2_W1(32'h3bfb0e7c), .K2_C2_W2(32'hbd3dc960), .K2_C2_W3(32'h3e268cd0), .K2_C2_W4(32'hbda64629), .K2_C2_W5(32'h3b2bfef2), .K2_C2_W6(32'hbe1734dc), .K2_C2_W7(32'hbe088c7f), .K2_C2_W8(32'h3dbd7743), 
		.K2_C3_W0(32'h3db7c4ce), .K2_C3_W1(32'hbdefb086), .K2_C3_W2(32'h3c72b89c), .K2_C3_W3(32'h3d9159a9), .K2_C3_W4(32'hbde8eb96), .K2_C3_W5(32'h3dd6ccb3), .K2_C3_W6(32'hbe1bf70e), .K2_C3_W7(32'hbda89052), .K2_C3_W8(32'hbdb7564b), 
		.K2_C4_W0(32'h3e1c5e13), .K2_C4_W1(32'h3d65bf7d), .K2_C4_W2(32'hbda4f891), .K2_C4_W3(32'h3d71e999), .K2_C4_W4(32'h3d3ed825), .K2_C4_W5(32'hbb3c3496), .K2_C4_W6(32'h3dbe40bf), .K2_C4_W7(32'h3d47a870), .K2_C4_W8(32'h3d7b8ca6), 
		.K2_C5_W0(32'hbe2e4e0a), .K2_C5_W1(32'hbd6b4fae), .K2_C5_W2(32'hbdf0b3ac), .K2_C5_W3(32'hbde8c7d6), .K2_C5_W4(32'hbdd2fba6), .K2_C5_W5(32'h3d47634d), .K2_C5_W6(32'h3d2ae2eb), .K2_C5_W7(32'hbda31aa9), .K2_C5_W8(32'hbdd242e6), 
		.K2_C6_W0(32'h3d12df27), .K2_C6_W1(32'hbdc96cc5), .K2_C6_W2(32'hbe132952), .K2_C6_W3(32'hbd66296a), .K2_C6_W4(32'hbda65ae3), .K2_C6_W5(32'h3de98f4f), .K2_C6_W6(32'hbdb93cd1), .K2_C6_W7(32'hbc62a671), .K2_C6_W8(32'hbc0f40d2), 
		.K2_C7_W0(32'hbd7503db), .K2_C7_W1(32'hbe094bea), .K2_C7_W2(32'h3d8fe39e), .K2_C7_W3(32'hbc939702), .K2_C7_W4(32'h3d2aa339), .K2_C7_W5(32'hbd89d5a7), .K2_C7_W6(32'hbe0b3368), .K2_C7_W7(32'hbe0aff2c), .K2_C7_W8(32'h3d3beba0), 
		.K2_C8_W0(32'hbce2d5c7), .K2_C8_W1(32'h3da3514f), .K2_C8_W2(32'hbc83c6d2), .K2_C8_W3(32'h3c77d052), .K2_C8_W4(32'h3d72d9a5), .K2_C8_W5(32'hbe017b4b), .K2_C8_W6(32'hbc9b49e1), .K2_C8_W7(32'h3da7facb), .K2_C8_W8(32'hbb2c6643), 
		.K2_C9_W0(32'hbde97907), .K2_C9_W1(32'hbc0ed706), .K2_C9_W2(32'hbc4e1f15), .K2_C9_W3(32'hbd4bf228), .K2_C9_W4(32'hbdda66b6), .K2_C9_W5(32'h3e053cfd), .K2_C9_W6(32'hbd8609f6), .K2_C9_W7(32'hbd9d567a), .K2_C9_W8(32'h3d825a40), 
		.K2_C10_W0(32'h3cf2b721), .K2_C10_W1(32'h3bf16a3e), .K2_C10_W2(32'h3d606535), .K2_C10_W3(32'h3e01d985), .K2_C10_W4(32'h3de2b414), .K2_C10_W5(32'hbdb3da14), .K2_C10_W6(32'hbdafb51e), .K2_C10_W7(32'h3d9ede76), .K2_C10_W8(32'h3cfa9286), 
		.K2_C11_W0(32'hbbc47771), .K2_C11_W1(32'h3e0b4690), .K2_C11_W2(32'h3de06121), .K2_C11_W3(32'h3c6a9ff2), .K2_C11_W4(32'h3d9b60f4), .K2_C11_W5(32'h3df73b1c), .K2_C11_W6(32'hbdd7ac3f), .K2_C11_W7(32'h3b85de2d), .K2_C11_W8(32'h3d952251), 
		.K2_C12_W0(32'h3d986fb9), .K2_C12_W1(32'h3da6c31c), .K2_C12_W2(32'hbca6c8e1), .K2_C12_W3(32'h3d48712c), .K2_C12_W4(32'h3d912c4d), .K2_C12_W5(32'hbd84e085), .K2_C12_W6(32'hbd42870a), .K2_C12_W7(32'hbc417437), .K2_C12_W8(32'h3c477a52), 
		.K2_C13_W0(32'h3d6a6202), .K2_C13_W1(32'hbe110da9), .K2_C13_W2(32'hbdf62631), .K2_C13_W3(32'hbde800fc), .K2_C13_W4(32'h3c600e2f), .K2_C13_W5(32'hbdd8b1c2), .K2_C13_W6(32'hbdc9e82d), .K2_C13_W7(32'hbd1d803b), .K2_C13_W8(32'h3d7de73c), 
		.K2_C14_W0(32'hbdf28df4), .K2_C14_W1(32'h3da7e4f7), .K2_C14_W2(32'hbddd7d9a), .K2_C14_W3(32'h3db5ba0b), .K2_C14_W4(32'h3e12f9ba), .K2_C14_W5(32'h3d5f4fe8), .K2_C14_W6(32'hbe12ce32), .K2_C14_W7(32'hbdca9a2c), .K2_C14_W8(32'h3cb8e5ad), 
		.K2_C15_W0(32'h3c37e1ec), .K2_C15_W1(32'h3e012fe0), .K2_C15_W2(32'h3e1bf461), .K2_C15_W3(32'h3e0cf3f1), .K2_C15_W4(32'hbced1be2), .K2_C15_W5(32'hbe20bcdf), .K2_C15_W6(32'h3df50600), .K2_C15_W7(32'hbccd6a82), .K2_C15_W8(32'hbda4c344), 
		.K2_BIAS (32'hbd11c529),

		.K3_C0_W0(32'h3de71966), .K3_C0_W1(32'h3c4e54c9), .K3_C0_W2(32'hbb200845), .K3_C0_W3(32'h3d14b66f), .K3_C0_W4(32'h3e008213), .K3_C0_W5(32'h3de0a198), .K3_C0_W6(32'hbe144726), .K3_C0_W7(32'h3de2cff1), .K3_C0_W8(32'hbd5264f8), 
		.K3_C1_W0(32'hbd03e19e), .K3_C1_W1(32'hbd7b3487), .K3_C1_W2(32'hbb9299b0), .K3_C1_W3(32'hbd812833), .K3_C1_W4(32'h3df631f7), .K3_C1_W5(32'hbd935a40), .K3_C1_W6(32'h3c6527ff), .K3_C1_W7(32'h3c958556), .K3_C1_W8(32'h3c489d0c), 
		.K3_C2_W0(32'hbdf25a68), .K3_C2_W1(32'hbcf8a739), .K3_C2_W2(32'h3dea2917), .K3_C2_W3(32'hbca0f332), .K3_C2_W4(32'h3c80b710), .K3_C2_W5(32'hbd983013), .K3_C2_W6(32'h3d967886), .K3_C2_W7(32'h3d1b1fcc), .K3_C2_W8(32'h3cd0765b), 
		.K3_C3_W0(32'h3d78c072), .K3_C3_W1(32'h3d75dc98), .K3_C3_W2(32'hbd8e59d3), .K3_C3_W3(32'h3dddedc6), .K3_C3_W4(32'hbe0cfcd2), .K3_C3_W5(32'h3dc3589b), .K3_C3_W6(32'h3e00c0f1), .K3_C3_W7(32'h3ca0629e), .K3_C3_W8(32'h3db9d850), 
		.K3_C4_W0(32'hbe0c492f), .K3_C4_W1(32'h3d0a1068), .K3_C4_W2(32'h3d175ab3), .K3_C4_W3(32'hbce1c9e2), .K3_C4_W4(32'h3e1d001e), .K3_C4_W5(32'h3aea4694), .K3_C4_W6(32'hbda80798), .K3_C4_W7(32'h3db4e52a), .K3_C4_W8(32'h3de9f5c9), 
		.K3_C5_W0(32'hbb487888), .K3_C5_W1(32'hbdd567dd), .K3_C5_W2(32'hbe217042), .K3_C5_W3(32'hbe4dfd6b), .K3_C5_W4(32'h3dc69121), .K3_C5_W5(32'hbc963c5d), .K3_C5_W6(32'hbe02a843), .K3_C5_W7(32'hbdb1964e), .K3_C5_W8(32'h3df9660d), 
		.K3_C6_W0(32'hbddc4284), .K3_C6_W1(32'h3d5f47c8), .K3_C6_W2(32'hbacfcf95), .K3_C6_W3(32'hbdcac846), .K3_C6_W4(32'hbdbbbbd3), .K3_C6_W5(32'hbd10c802), .K3_C6_W6(32'hbd97a721), .K3_C6_W7(32'hbd86a943), .K3_C6_W8(32'h3ddc49f6), 
		.K3_C7_W0(32'h3da1f76d), .K3_C7_W1(32'h3db6e7db), .K3_C7_W2(32'hbd9400f0), .K3_C7_W3(32'hbd91f388), .K3_C7_W4(32'hbd5fd51f), .K3_C7_W5(32'h3db7039a), .K3_C7_W6(32'hbdfc147e), .K3_C7_W7(32'h3d4114f7), .K3_C7_W8(32'hbd77d8b8), 
		.K3_C8_W0(32'hbd8b5531), .K3_C8_W1(32'h3d9192c2), .K3_C8_W2(32'hbde4875c), .K3_C8_W3(32'h3dcc229a), .K3_C8_W4(32'h3c44e486), .K3_C8_W5(32'h3dd0a01a), .K3_C8_W6(32'h3ddb38d5), .K3_C8_W7(32'hbd2c9d79), .K3_C8_W8(32'hbd5497ce), 
		.K3_C9_W0(32'hbdefb227), .K3_C9_W1(32'hbb28e33f), .K3_C9_W2(32'hbdc0bd04), .K3_C9_W3(32'hbdf7a228), .K3_C9_W4(32'h3ddf64f4), .K3_C9_W5(32'h3d50741d), .K3_C9_W6(32'hbe09949f), .K3_C9_W7(32'hbce08f1d), .K3_C9_W8(32'h3e0f0c0f), 
		.K3_C10_W0(32'h3d8c842c), .K3_C10_W1(32'h3e0cebdd), .K3_C10_W2(32'hbdfde30d), .K3_C10_W3(32'h3ca29213), .K3_C10_W4(32'hbe14ab77), .K3_C10_W5(32'hbd9626b1), .K3_C10_W6(32'hbd6fc79e), .K3_C10_W7(32'h3d94ba85), .K3_C10_W8(32'hbddaa7e7), 
		.K3_C11_W0(32'h3e025c7f), .K3_C11_W1(32'h3e11cf34), .K3_C11_W2(32'hbcbdbf6c), .K3_C11_W3(32'h3bebe990), .K3_C11_W4(32'h3db59929), .K3_C11_W5(32'hbdb55df5), .K3_C11_W6(32'h3dd189ed), .K3_C11_W7(32'h3c645877), .K3_C11_W8(32'h3b17a42b), 
		.K3_C12_W0(32'h3d6fa46e), .K3_C12_W1(32'h3dae1890), .K3_C12_W2(32'hbdb1bf9d), .K3_C12_W3(32'h3cfe2a05), .K3_C12_W4(32'h3dc23ee6), .K3_C12_W5(32'h3c2ddfc8), .K3_C12_W6(32'hbe0de6ca), .K3_C12_W7(32'hbc3f0187), .K3_C12_W8(32'h3d6b6963), 
		.K3_C13_W0(32'hbd937f0b), .K3_C13_W1(32'hbcd15af3), .K3_C13_W2(32'hbca6d011), .K3_C13_W3(32'h3ddd8274), .K3_C13_W4(32'hbdc836fb), .K3_C13_W5(32'hbe08fb5c), .K3_C13_W6(32'h3ddc5396), .K3_C13_W7(32'hbbef6939), .K3_C13_W8(32'h3d12ccbf), 
		.K3_C14_W0(32'h3d74485d), .K3_C14_W1(32'h3e0bcd83), .K3_C14_W2(32'h3da3cb57), .K3_C14_W3(32'hbe121b77), .K3_C14_W4(32'hbdaabb83), .K3_C14_W5(32'h3d8f9362), .K3_C14_W6(32'h3dcdf994), .K3_C14_W7(32'h3df579d9), .K3_C14_W8(32'h3ddbdead), 
		.K3_C15_W0(32'hbd345122), .K3_C15_W1(32'hbc81785d), .K3_C15_W2(32'hbe010d6d), .K3_C15_W3(32'h3d9ae5df), .K3_C15_W4(32'h3de05984), .K3_C15_W5(32'hbd8ba64e), .K3_C15_W6(32'hbd4333ae), .K3_C15_W7(32'h3d9a7ccd), .K3_C15_W8(32'h3d8fc3b7), 
		.K3_BIAS (32'hbd30d3d2),

		.K4_C0_W0(32'hbe08ade2), .K4_C0_W1(32'h3d7df7f2), .K4_C0_W2(32'hbe0d3410), .K4_C0_W3(32'h3d048b16), .K4_C0_W4(32'h3d527c5c), .K4_C0_W5(32'hbde982f3), .K4_C0_W6(32'hb9ebf0c5), .K4_C0_W7(32'h3d4f4a83), .K4_C0_W8(32'hbcac41a8), 
		.K4_C1_W0(32'h3b15d3be), .K4_C1_W1(32'hbe0abc1a), .K4_C1_W2(32'h3c55e871), .K4_C1_W3(32'hbcaf2386), .K4_C1_W4(32'h3dc140a4), .K4_C1_W5(32'hbde57c4d), .K4_C1_W6(32'hbbb176bc), .K4_C1_W7(32'h3db2a526), .K4_C1_W8(32'h3c31f5e8), 
		.K4_C2_W0(32'hbd54334e), .K4_C2_W1(32'h3b998466), .K4_C2_W2(32'hbd342466), .K4_C2_W3(32'h3e32a92c), .K4_C2_W4(32'hbd14e984), .K4_C2_W5(32'hbdb11c20), .K4_C2_W6(32'hbd8b9626), .K4_C2_W7(32'h3dac886a), .K4_C2_W8(32'h3cc75bf2), 
		.K4_C3_W0(32'h3dc96ad6), .K4_C3_W1(32'h3c9b98e1), .K4_C3_W2(32'hbe07ca6d), .K4_C3_W3(32'hbd0188bc), .K4_C3_W4(32'hbd1ec18b), .K4_C3_W5(32'hbca2dea7), .K4_C3_W6(32'hbdbc9ac2), .K4_C3_W7(32'hbbd726b0), .K4_C3_W8(32'hbdfd252f), 
		.K4_C4_W0(32'hbdaf0f57), .K4_C4_W1(32'h3d94088f), .K4_C4_W2(32'h3e1c3c1e), .K4_C4_W3(32'h3cce8eb2), .K4_C4_W4(32'hbe09d416), .K4_C4_W5(32'hbd8dc10a), .K4_C4_W6(32'h3d3388f1), .K4_C4_W7(32'h3d73724c), .K4_C4_W8(32'hbdcb3ad2), 
		.K4_C5_W0(32'hbd971f7e), .K4_C5_W1(32'h3d4aaa38), .K4_C5_W2(32'hbdb65812), .K4_C5_W3(32'hbd17da72), .K4_C5_W4(32'hbd17363f), .K4_C5_W5(32'h3dd4fab8), .K4_C5_W6(32'h3cfaac79), .K4_C5_W7(32'hbda1ccde), .K4_C5_W8(32'hbca74510), 
		.K4_C6_W0(32'hbdce9e19), .K4_C6_W1(32'h3df0e38c), .K4_C6_W2(32'h3c1799ec), .K4_C6_W3(32'hbd1403b3), .K4_C6_W4(32'hbd293f85), .K4_C6_W5(32'h3dc85ee7), .K4_C6_W6(32'hbd36db78), .K4_C6_W7(32'h3e12f089), .K4_C6_W8(32'hbd4a5d8d), 
		.K4_C7_W0(32'hbca38708), .K4_C7_W1(32'h3c964902), .K4_C7_W2(32'h3dd978d7), .K4_C7_W3(32'h3d258883), .K4_C7_W4(32'h3b1510e5), .K4_C7_W5(32'h3d05e81e), .K4_C7_W6(32'hbd2d214b), .K4_C7_W7(32'h3d7365d6), .K4_C7_W8(32'hbb91faf8), 
		.K4_C8_W0(32'hbda81680), .K4_C8_W1(32'h3d271e50), .K4_C8_W2(32'hbd75b5a0), .K4_C8_W3(32'hbd884596), .K4_C8_W4(32'h3d3b1c54), .K4_C8_W5(32'h3e030bdf), .K4_C8_W6(32'h3b50c0d0), .K4_C8_W7(32'h3d0d918a), .K4_C8_W8(32'hbd5a8127), 
		.K4_C9_W0(32'h3dbdd780), .K4_C9_W1(32'hbdf37374), .K4_C9_W2(32'h3c8006e7), .K4_C9_W3(32'hbd9f2563), .K4_C9_W4(32'h3d2c13a7), .K4_C9_W5(32'h3db207dd), .K4_C9_W6(32'h3e1715c3), .K4_C9_W7(32'h3e30e42f), .K4_C9_W8(32'h3df74165), 
		.K4_C10_W0(32'h3ddd3342), .K4_C10_W1(32'h3d908132), .K4_C10_W2(32'hbe106f42), .K4_C10_W3(32'h3df33c47), .K4_C10_W4(32'hbda3fac8), .K4_C10_W5(32'hbd0fea60), .K4_C10_W6(32'hbdd91451), .K4_C10_W7(32'hbc860eb7), .K4_C10_W8(32'hbda55ea2), 
		.K4_C11_W0(32'h3de47e5a), .K4_C11_W1(32'hbdd4038a), .K4_C11_W2(32'hbdd56bfe), .K4_C11_W3(32'hbd51dac1), .K4_C11_W4(32'h3daac608), .K4_C11_W5(32'h3c41c049), .K4_C11_W6(32'hbe01c50d), .K4_C11_W7(32'hbb0cb4a2), .K4_C11_W8(32'hbdd0e1a9), 
		.K4_C12_W0(32'hbe09f545), .K4_C12_W1(32'h3e001e79), .K4_C12_W2(32'hbbf76e21), .K4_C12_W3(32'hbd4712fc), .K4_C12_W4(32'hbe05090d), .K4_C12_W5(32'h3dbee7b2), .K4_C12_W6(32'h3dae0beb), .K4_C12_W7(32'hbd6422e6), .K4_C12_W8(32'h3cea01b0), 
		.K4_C13_W0(32'hbccd6e70), .K4_C13_W1(32'hbdd8c3a1), .K4_C13_W2(32'hbdb42a8e), .K4_C13_W3(32'h3de0f6a5), .K4_C13_W4(32'hbe20f047), .K4_C13_W5(32'hbe0c16e6), .K4_C13_W6(32'hbddf9cde), .K4_C13_W7(32'hbe08a6b0), .K4_C13_W8(32'h3e0e62a8), 
		.K4_C14_W0(32'h3dac62ea), .K4_C14_W1(32'h3d8f2664), .K4_C14_W2(32'h3b1b2b27), .K4_C14_W3(32'h3cdaf1f9), .K4_C14_W4(32'h3dbb036e), .K4_C14_W5(32'hbdbbc1f5), .K4_C14_W6(32'hbdac8b74), .K4_C14_W7(32'h3d74e3dd), .K4_C14_W8(32'h3d04e637), 
		.K4_C15_W0(32'hbc9185c0), .K4_C15_W1(32'hbe14dd19), .K4_C15_W2(32'hbcd5b0b1), .K4_C15_W3(32'h3e0a2cbb), .K4_C15_W4(32'h3da0da03), .K4_C15_W5(32'h3dae33a0), .K4_C15_W6(32'hbdcfcb62), .K4_C15_W7(32'hbc170599), .K4_C15_W8(32'h3d87cba4), 
		.K4_BIAS (32'h3d23b5d8),

		.K5_C0_W0(32'h3c3f10bc), .K5_C0_W1(32'h3e14e232), .K5_C0_W2(32'h3db0c696), .K5_C0_W3(32'h3e26d929), .K5_C0_W4(32'h3d80dd6c), .K5_C0_W5(32'h3e2fc3bd), .K5_C0_W6(32'h3e2f82c5), .K5_C0_W7(32'hbd815184), .K5_C0_W8(32'h3cd9f59a), 
		.K5_C1_W0(32'hbe0b57af), .K5_C1_W1(32'h3de531f3), .K5_C1_W2(32'h3dec77f2), .K5_C1_W3(32'h3c0d87d4), .K5_C1_W4(32'h3cf61733), .K5_C1_W5(32'hbdad6f0e), .K5_C1_W6(32'h3dfec6ac), .K5_C1_W7(32'hbd9e422a), .K5_C1_W8(32'h3d285d1d), 
		.K5_C2_W0(32'h3d9968e6), .K5_C2_W1(32'h3bd4c98f), .K5_C2_W2(32'hbd0b7788), .K5_C2_W3(32'h3c55fe52), .K5_C2_W4(32'h3c9bc008), .K5_C2_W5(32'h3d6229b3), .K5_C2_W6(32'hbcbb0a18), .K5_C2_W7(32'h3dcab95d), .K5_C2_W8(32'hbd598fd4), 
		.K5_C3_W0(32'hbdd6c5d5), .K5_C3_W1(32'hbd1926bb), .K5_C3_W2(32'hbd5542ec), .K5_C3_W3(32'hbdd1fd4d), .K5_C3_W4(32'hbd66e33d), .K5_C3_W5(32'h3d497704), .K5_C3_W6(32'hbcc50630), .K5_C3_W7(32'hbe1a68a1), .K5_C3_W8(32'h3dc45e76), 
		.K5_C4_W0(32'hbd0e37d9), .K5_C4_W1(32'h3e20c842), .K5_C4_W2(32'hbd470aba), .K5_C4_W3(32'hbd873588), .K5_C4_W4(32'hbc980314), .K5_C4_W5(32'h3c184a4a), .K5_C4_W6(32'h3d4c5b22), .K5_C4_W7(32'hbdf80bb3), .K5_C4_W8(32'hbe02b40d), 
		.K5_C5_W0(32'hbdb81b0f), .K5_C5_W1(32'hbd9adee1), .K5_C5_W2(32'h3ddc7c7a), .K5_C5_W3(32'hbd94fc11), .K5_C5_W4(32'hbd09f6ef), .K5_C5_W5(32'h3db58e8a), .K5_C5_W6(32'hbdcd78ae), .K5_C5_W7(32'h3d61578d), .K5_C5_W8(32'hbb8bcb00), 
		.K5_C6_W0(32'hbc26513f), .K5_C6_W1(32'hbd90eeb5), .K5_C6_W2(32'hbd2dfae0), .K5_C6_W3(32'hbc7a3396), .K5_C6_W4(32'h3e03bccb), .K5_C6_W5(32'hbc68232d), .K5_C6_W6(32'hbda53874), .K5_C6_W7(32'h3d7ccc73), .K5_C6_W8(32'hbdf78434), 
		.K5_C7_W0(32'h3b3f1328), .K5_C7_W1(32'hbc974ff2), .K5_C7_W2(32'h3d770b81), .K5_C7_W3(32'hbc2ff856), .K5_C7_W4(32'hbdffcf9a), .K5_C7_W5(32'h3de470ac), .K5_C7_W6(32'hbe0bf31c), .K5_C7_W7(32'h3d7fb742), .K5_C7_W8(32'hbdadb4a4), 
		.K5_C8_W0(32'hbdfe99e1), .K5_C8_W1(32'hbd97d343), .K5_C8_W2(32'hbd303dc6), .K5_C8_W3(32'hbe27c3b7), .K5_C8_W4(32'hbda84036), .K5_C8_W5(32'hbdd4224d), .K5_C8_W6(32'h3cf5ea33), .K5_C8_W7(32'hbe2964f9), .K5_C8_W8(32'hbd6f0e10), 
		.K5_C9_W0(32'h3d730d95), .K5_C9_W1(32'hbd9c2a57), .K5_C9_W2(32'hbd1f6781), .K5_C9_W3(32'h3c922e0a), .K5_C9_W4(32'h3d5f73a0), .K5_C9_W5(32'hbd186756), .K5_C9_W6(32'h3c733e75), .K5_C9_W7(32'h3e187bca), .K5_C9_W8(32'h3e02a414), 
		.K5_C10_W0(32'hbd51396c), .K5_C10_W1(32'h3e06c691), .K5_C10_W2(32'h3d8d3553), .K5_C10_W3(32'h3dd627ce), .K5_C10_W4(32'hbda78f4c), .K5_C10_W5(32'hbd0c7858), .K5_C10_W6(32'hbe02ed78), .K5_C10_W7(32'hbd85a871), .K5_C10_W8(32'hbe175c6b), 
		.K5_C11_W0(32'h3d8e3ab0), .K5_C11_W1(32'hbe0b0352), .K5_C11_W2(32'hbdc5ebeb), .K5_C11_W3(32'hbc8c624b), .K5_C11_W4(32'hbdf27ad0), .K5_C11_W5(32'hbdd5c527), .K5_C11_W6(32'h3ca79768), .K5_C11_W7(32'hbda8e369), .K5_C11_W8(32'hbd522d2c), 
		.K5_C12_W0(32'hbcd431dc), .K5_C12_W1(32'hbdd4ed82), .K5_C12_W2(32'h3d8e068c), .K5_C12_W3(32'hbdb64bfb), .K5_C12_W4(32'h3df0674f), .K5_C12_W5(32'h3cb44dec), .K5_C12_W6(32'h3d03e5e3), .K5_C12_W7(32'h3da4802e), .K5_C12_W8(32'h3d893ab6), 
		.K5_C13_W0(32'hbc41fae6), .K5_C13_W1(32'h3df1af7b), .K5_C13_W2(32'h3dd0acbc), .K5_C13_W3(32'hbc809aae), .K5_C13_W4(32'hbc6ec45d), .K5_C13_W5(32'hbc37cc9f), .K5_C13_W6(32'hbbfb7843), .K5_C13_W7(32'hbdb35744), .K5_C13_W8(32'hbdc6468b), 
		.K5_C14_W0(32'h3de3e923), .K5_C14_W1(32'hbdd27301), .K5_C14_W2(32'h3d6e1e70), .K5_C14_W3(32'hbd215492), .K5_C14_W4(32'hbd63c3dd), .K5_C14_W5(32'h3bb223fd), .K5_C14_W6(32'h3d94ac38), .K5_C14_W7(32'hbb19fbeb), .K5_C14_W8(32'hbdb01cf3), 
		.K5_C15_W0(32'hbdd32bf4), .K5_C15_W1(32'hbd4ac41e), .K5_C15_W2(32'hbd81c730), .K5_C15_W3(32'h3c2cad43), .K5_C15_W4(32'h3d53716e), .K5_C15_W5(32'hbd2316de), .K5_C15_W6(32'hbdf923d6), .K5_C15_W7(32'h3bfe14ed), .K5_C15_W8(32'hbd7cc74a), 
		.K5_BIAS (32'hbcc1bc3e),

		.K6_C0_W0(32'hbdeaac23), .K6_C0_W1(32'h3cbcbd65), .K6_C0_W2(32'h3d413e37), .K6_C0_W3(32'hbdcd0db7), .K6_C0_W4(32'hbd8992ca), .K6_C0_W5(32'h3d0f5418), .K6_C0_W6(32'h3cdea13b), .K6_C0_W7(32'h3dce5d23), .K6_C0_W8(32'hbcf8e580), 
		.K6_C1_W0(32'h3dffc004), .K6_C1_W1(32'h3e11d505), .K6_C1_W2(32'h3dcf54a8), .K6_C1_W3(32'h3cbc5d41), .K6_C1_W4(32'hbd81a468), .K6_C1_W5(32'hbd7c7ee6), .K6_C1_W6(32'hbce09e07), .K6_C1_W7(32'hbdcdc4bb), .K6_C1_W8(32'hbd6d8007), 
		.K6_C2_W0(32'h3d8108dc), .K6_C2_W1(32'h3dcca3ca), .K6_C2_W2(32'h3deb45cb), .K6_C2_W3(32'h3d4d5de6), .K6_C2_W4(32'hbda91172), .K6_C2_W5(32'hbded6264), .K6_C2_W6(32'hbdc0d0d7), .K6_C2_W7(32'hbdcff946), .K6_C2_W8(32'hbcd58a7c), 
		.K6_C3_W0(32'hbceedc59), .K6_C3_W1(32'hbde576ac), .K6_C3_W2(32'hbc0cfe27), .K6_C3_W3(32'h3e022a87), .K6_C3_W4(32'hbd306b48), .K6_C3_W5(32'h3e014ba6), .K6_C3_W6(32'hbce98b04), .K6_C3_W7(32'h3d5682fd), .K6_C3_W8(32'hbd99f5dc), 
		.K6_C4_W0(32'h3d6a9f9c), .K6_C4_W1(32'h3c0810b8), .K6_C4_W2(32'hbd2a0dbf), .K6_C4_W3(32'hbd8475bf), .K6_C4_W4(32'hbe0b0b58), .K6_C4_W5(32'hbd83e9a8), .K6_C4_W6(32'h3cd73a38), .K6_C4_W7(32'hbe003cdf), .K6_C4_W8(32'h3cf4cf17), 
		.K6_C5_W0(32'hbddc5508), .K6_C5_W1(32'hbe2a5d71), .K6_C5_W2(32'h3cbd7300), .K6_C5_W3(32'hbc1754f8), .K6_C5_W4(32'hbe1b09d7), .K6_C5_W5(32'hbd2705b7), .K6_C5_W6(32'hbd45d01b), .K6_C5_W7(32'hbe1024ac), .K6_C5_W8(32'hbe2353d5), 
		.K6_C6_W0(32'hbdaace9b), .K6_C6_W1(32'h3e07b2d5), .K6_C6_W2(32'hbd8a888d), .K6_C6_W3(32'h3cd389fb), .K6_C6_W4(32'h3c6eef00), .K6_C6_W5(32'h3ddfa0ef), .K6_C6_W6(32'h3c09d199), .K6_C6_W7(32'h3e167069), .K6_C6_W8(32'h3d026410), 
		.K6_C7_W0(32'hbdfed26b), .K6_C7_W1(32'hbd7e05a1), .K6_C7_W2(32'hbe043fea), .K6_C7_W3(32'h3e138f7e), .K6_C7_W4(32'hbd9ef7b9), .K6_C7_W5(32'hbd9b3ba9), .K6_C7_W6(32'h3db803f2), .K6_C7_W7(32'h3e059e4e), .K6_C7_W8(32'h3d461777), 
		.K6_C8_W0(32'h3dcf9fb3), .K6_C8_W1(32'hbc5b1c8c), .K6_C8_W2(32'hbd91be69), .K6_C8_W3(32'h3d9a17de), .K6_C8_W4(32'hbdd8ce0f), .K6_C8_W5(32'h3d9ad010), .K6_C8_W6(32'h3e1cb683), .K6_C8_W7(32'h3c4993ea), .K6_C8_W8(32'h3d1a521d), 
		.K6_C9_W0(32'hbd0b1e0f), .K6_C9_W1(32'hbc93313d), .K6_C9_W2(32'hbe0297d0), .K6_C9_W3(32'h3e1713ed), .K6_C9_W4(32'h3e176213), .K6_C9_W5(32'h3c20485d), .K6_C9_W6(32'h3e13ff5c), .K6_C9_W7(32'h3d677bcf), .K6_C9_W8(32'h3d49a2c3), 
		.K6_C10_W0(32'h3db16d97), .K6_C10_W1(32'h3cdc8118), .K6_C10_W2(32'hbdac3a71), .K6_C10_W3(32'h3dfcf107), .K6_C10_W4(32'hbde03133), .K6_C10_W5(32'hbc7feb93), .K6_C10_W6(32'hbde6c39b), .K6_C10_W7(32'hbd0acfb0), .K6_C10_W8(32'hbd029172), 
		.K6_C11_W0(32'h3d0efecd), .K6_C11_W1(32'h3d5e9b84), .K6_C11_W2(32'h3ded985d), .K6_C11_W3(32'h3c2538d9), .K6_C11_W4(32'h3e05c025), .K6_C11_W5(32'hbd3c0918), .K6_C11_W6(32'hbd980d6a), .K6_C11_W7(32'h3e109981), .K6_C11_W8(32'hbe059039), 
		.K6_C12_W0(32'hbe0d9b70), .K6_C12_W1(32'hbe06811b), .K6_C12_W2(32'h3dcb8cde), .K6_C12_W3(32'hbc9ff027), .K6_C12_W4(32'h3e00ee70), .K6_C12_W5(32'h3dfd8519), .K6_C12_W6(32'hbc3ce3e2), .K6_C12_W7(32'h3be72d1f), .K6_C12_W8(32'hbb89a982), 
		.K6_C13_W0(32'hbd0a1513), .K6_C13_W1(32'h3d39a140), .K6_C13_W2(32'hbd1aa89c), .K6_C13_W3(32'hbd4b452d), .K6_C13_W4(32'hbca83244), .K6_C13_W5(32'hbd63ef59), .K6_C13_W6(32'hbdf60a9f), .K6_C13_W7(32'h3af49e06), .K6_C13_W8(32'h3e0b10aa), 
		.K6_C14_W0(32'h3c143138), .K6_C14_W1(32'hbe18e50e), .K6_C14_W2(32'hbd9764f0), .K6_C14_W3(32'h3da5354a), .K6_C14_W4(32'h3d5ad566), .K6_C14_W5(32'hbd8ea386), .K6_C14_W6(32'hbcaf4b28), .K6_C14_W7(32'h3d0e9d18), .K6_C14_W8(32'h3dc4a734), 
		.K6_C15_W0(32'hbe0bb494), .K6_C15_W1(32'h3d42eaf0), .K6_C15_W2(32'h3c8f796f), .K6_C15_W3(32'h3c050038), .K6_C15_W4(32'hbb98601e), .K6_C15_W5(32'hbe0dd7e4), .K6_C15_W6(32'hbd52899c), .K6_C15_W7(32'h3d4d6ed3), .K6_C15_W8(32'hbd7d35c6), 
		.K6_BIAS (32'h3c139d17),

		.K7_C0_W0(32'h3d9f3baa), .K7_C0_W1(32'h3de0fccf), .K7_C0_W2(32'h3d3d520f), .K7_C0_W3(32'h3de453e6), .K7_C0_W4(32'h3dce258d), .K7_C0_W5(32'hbdf49198), .K7_C0_W6(32'h3df13229), .K7_C0_W7(32'h3d74b89e), .K7_C0_W8(32'hbdc77495), 
		.K7_C1_W0(32'h3d87dd9d), .K7_C1_W1(32'hbdb1603c), .K7_C1_W2(32'hbdcff5a8), .K7_C1_W3(32'hbdb3bf18), .K7_C1_W4(32'h3cbe1857), .K7_C1_W5(32'h3d66f0c7), .K7_C1_W6(32'h3d33197a), .K7_C1_W7(32'h3de12d9a), .K7_C1_W8(32'hbc9755aa), 
		.K7_C2_W0(32'hbcee2b78), .K7_C2_W1(32'h3e14af2a), .K7_C2_W2(32'h3d4e56a1), .K7_C2_W3(32'hbdab1f41), .K7_C2_W4(32'h3da216be), .K7_C2_W5(32'h3dfe37e7), .K7_C2_W6(32'h3befa107), .K7_C2_W7(32'h3dfc6aca), .K7_C2_W8(32'h3dcd8edd), 
		.K7_C3_W0(32'h3bd980d6), .K7_C3_W1(32'hbd347827), .K7_C3_W2(32'h3d41516c), .K7_C3_W3(32'h3d5814dd), .K7_C3_W4(32'h3e1c3cb5), .K7_C3_W5(32'hbd87b4a8), .K7_C3_W6(32'h3c9e057b), .K7_C3_W7(32'hbde2ae6f), .K7_C3_W8(32'hbc91c630), 
		.K7_C4_W0(32'h3defb562), .K7_C4_W1(32'h3c6b3c9c), .K7_C4_W2(32'hbde2b5f6), .K7_C4_W3(32'hbd8130dc), .K7_C4_W4(32'hbe18924f), .K7_C4_W5(32'h3a50765b), .K7_C4_W6(32'h3c1a0d32), .K7_C4_W7(32'hbd8db15b), .K7_C4_W8(32'hbdba8c36), 
		.K7_C5_W0(32'h3df59dbe), .K7_C5_W1(32'hbe096f55), .K7_C5_W2(32'hbe0f4ea8), .K7_C5_W3(32'hbdc6894d), .K7_C5_W4(32'hbce5bba3), .K7_C5_W5(32'hbd8af31d), .K7_C5_W6(32'hbdd748d5), .K7_C5_W7(32'h3e0ca7bc), .K7_C5_W8(32'hbc9c2b95), 
		.K7_C6_W0(32'hbe0883b3), .K7_C6_W1(32'h3c9668b1), .K7_C6_W2(32'h3d6456dc), .K7_C6_W3(32'hbdb72fdc), .K7_C6_W4(32'h3cf15790), .K7_C6_W5(32'h3bfb984d), .K7_C6_W6(32'h3caafe4a), .K7_C6_W7(32'h3b363904), .K7_C6_W8(32'h3dad507b), 
		.K7_C7_W0(32'h3dfd2fdf), .K7_C7_W1(32'hbd8fd408), .K7_C7_W2(32'hbde0d670), .K7_C7_W3(32'hbdca8c49), .K7_C7_W4(32'h3df19729), .K7_C7_W5(32'h3d1e5b44), .K7_C7_W6(32'hbbc7f49e), .K7_C7_W7(32'h3c737c75), .K7_C7_W8(32'hbe00c9fc), 
		.K7_C8_W0(32'hbb32c679), .K7_C8_W1(32'h3d31581c), .K7_C8_W2(32'hbda06fe0), .K7_C8_W3(32'hbe11d63e), .K7_C8_W4(32'hbcf7b21a), .K7_C8_W5(32'hbdfaac61), .K7_C8_W6(32'hbe0b1327), .K7_C8_W7(32'h3ddb2ff3), .K7_C8_W8(32'hbde60240), 
		.K7_C9_W0(32'hbe1c80f1), .K7_C9_W1(32'h3bd50168), .K7_C9_W2(32'h3d12351b), .K7_C9_W3(32'h3b24cdd5), .K7_C9_W4(32'hbd560615), .K7_C9_W5(32'hbe12d342), .K7_C9_W6(32'h3ccb0896), .K7_C9_W7(32'h3de73926), .K7_C9_W8(32'hbdee5c4b), 
		.K7_C10_W0(32'h3d2f6546), .K7_C10_W1(32'h3bf53b61), .K7_C10_W2(32'h3d939e68), .K7_C10_W3(32'hbdcbf99a), .K7_C10_W4(32'h3d9dd4ac), .K7_C10_W5(32'h3d95a17d), .K7_C10_W6(32'h3dbf2468), .K7_C10_W7(32'hbc921dcf), .K7_C10_W8(32'h3d877ba0), 
		.K7_C11_W0(32'hbd40a3d7), .K7_C11_W1(32'h3da73015), .K7_C11_W2(32'hbda51564), .K7_C11_W3(32'h3df29502), .K7_C11_W4(32'h3da91749), .K7_C11_W5(32'h3de98a1e), .K7_C11_W6(32'hbd99411f), .K7_C11_W7(32'hbc8f88eb), .K7_C11_W8(32'hbce5e45d), 
		.K7_C12_W0(32'h3c13a990), .K7_C12_W1(32'hbdbe2e6d), .K7_C12_W2(32'hbe21fb20), .K7_C12_W3(32'hbd7f47cc), .K7_C12_W4(32'hbe0e71b9), .K7_C12_W5(32'hbdd5c3bd), .K7_C12_W6(32'hbd6d3f4a), .K7_C12_W7(32'hbdd833c9), .K7_C12_W8(32'h3dbde849), 
		.K7_C13_W0(32'hbd110fb3), .K7_C13_W1(32'hbe159e93), .K7_C13_W2(32'hbdc8bd3c), .K7_C13_W3(32'hbe17e8a5), .K7_C13_W4(32'hbe21c0ef), .K7_C13_W5(32'h3c5ad325), .K7_C13_W6(32'hbdb8fb30), .K7_C13_W7(32'hbe18889f), .K7_C13_W8(32'hbe01887e), 
		.K7_C14_W0(32'h3d1005b7), .K7_C14_W1(32'h3e031976), .K7_C14_W2(32'hbcc70ed3), .K7_C14_W3(32'hbc8f5334), .K7_C14_W4(32'hbd90bb35), .K7_C14_W5(32'h3e12218f), .K7_C14_W6(32'h3d9a3f17), .K7_C14_W7(32'hbe1c4cea), .K7_C14_W8(32'h3d29b8b3), 
		.K7_C15_W0(32'h3de24c4d), .K7_C15_W1(32'hbd8535af), .K7_C15_W2(32'h3db04e29), .K7_C15_W3(32'h3ce2c676), .K7_C15_W4(32'hbd8e4a58), .K7_C15_W5(32'hbd07cbf0), .K7_C15_W6(32'h3cf309ed), .K7_C15_W7(32'h3d036b5e), .K7_C15_W8(32'hbc18f7bd), 
		.K7_BIAS (32'hbaa82ac9),

		.K8_C0_W0(32'h3dbd6642), .K8_C0_W1(32'h3ca94a00), .K8_C0_W2(32'hbdadddc3), .K8_C0_W3(32'hbd48e2c8), .K8_C0_W4(32'hbcf39be8), .K8_C0_W5(32'hbd43a1e9), .K8_C0_W6(32'hbd1846e2), .K8_C0_W7(32'h3e0943b2), .K8_C0_W8(32'h3d9bc349), 
		.K8_C1_W0(32'h3dab8472), .K8_C1_W1(32'h3e09f0b8), .K8_C1_W2(32'hbdf87a0f), .K8_C1_W3(32'hbde9ec2f), .K8_C1_W4(32'h3c85f2e5), .K8_C1_W5(32'hba2c9c3a), .K8_C1_W6(32'hbc42a9a5), .K8_C1_W7(32'h3e062a61), .K8_C1_W8(32'h3e062c1c), 
		.K8_C2_W0(32'h3d9f7a23), .K8_C2_W1(32'hbdfe5fbc), .K8_C2_W2(32'hbdd649c3), .K8_C2_W3(32'h3d324c6c), .K8_C2_W4(32'h3e0fe1bc), .K8_C2_W5(32'hbe041386), .K8_C2_W6(32'h3d7096b0), .K8_C2_W7(32'h3cffde47), .K8_C2_W8(32'h3e04005a), 
		.K8_C3_W0(32'hbd07f75f), .K8_C3_W1(32'h3dc9ebfb), .K8_C3_W2(32'h3d7593bf), .K8_C3_W3(32'h3dba560a), .K8_C3_W4(32'h3ca180ca), .K8_C3_W5(32'h3da12882), .K8_C3_W6(32'h3d675ae7), .K8_C3_W7(32'hbd901dba), .K8_C3_W8(32'hbdaa52b5), 
		.K8_C4_W0(32'hbd824d1e), .K8_C4_W1(32'hbd224ea6), .K8_C4_W2(32'h3e25955a), .K8_C4_W3(32'hbd3e3116), .K8_C4_W4(32'hbdbd4d83), .K8_C4_W5(32'hbda7f0b6), .K8_C4_W6(32'h3de72f43), .K8_C4_W7(32'h3e0f73b0), .K8_C4_W8(32'hbde1fda8), 
		.K8_C5_W0(32'h3df04676), .K8_C5_W1(32'h3d3a3a23), .K8_C5_W2(32'h3c82d870), .K8_C5_W3(32'hbd943b28), .K8_C5_W4(32'h3d3ce2b1), .K8_C5_W5(32'hbe04fae9), .K8_C5_W6(32'h3db53c6a), .K8_C5_W7(32'h3cbdcf03), .K8_C5_W8(32'h3dd7323a), 
		.K8_C6_W0(32'h3dd59c42), .K8_C6_W1(32'h3dc570c1), .K8_C6_W2(32'hbcc5c297), .K8_C6_W3(32'hbda84223), .K8_C6_W4(32'hbde2894d), .K8_C6_W5(32'h3e1289b6), .K8_C6_W6(32'hbda0fb80), .K8_C6_W7(32'hbe0261b7), .K8_C6_W8(32'hbca6063e), 
		.K8_C7_W0(32'hbda632d4), .K8_C7_W1(32'h3d1d740c), .K8_C7_W2(32'hbbf82ef3), .K8_C7_W3(32'hbda621b5), .K8_C7_W4(32'hbd9ccac2), .K8_C7_W5(32'hbc8b1664), .K8_C7_W6(32'h3dca5aad), .K8_C7_W7(32'h3d3efe3d), .K8_C7_W8(32'h3dde66b0), 
		.K8_C8_W0(32'hbd829f64), .K8_C8_W1(32'h3d29a686), .K8_C8_W2(32'h3e195524), .K8_C8_W3(32'h3cdf2adc), .K8_C8_W4(32'h3e0d09b0), .K8_C8_W5(32'hbdf7733f), .K8_C8_W6(32'hbd222694), .K8_C8_W7(32'hbdb799ec), .K8_C8_W8(32'hbd930e78), 
		.K8_C9_W0(32'h3d128032), .K8_C9_W1(32'h3da38857), .K8_C9_W2(32'hbe069963), .K8_C9_W3(32'hbc56b70b), .K8_C9_W4(32'hbdad0a5e), .K8_C9_W5(32'hbe17fc59), .K8_C9_W6(32'hbe2be754), .K8_C9_W7(32'h3c07d9fe), .K8_C9_W8(32'hbc8de9d1), 
		.K8_C10_W0(32'hbce9c349), .K8_C10_W1(32'hbda58915), .K8_C10_W2(32'h3dbdebb8), .K8_C10_W3(32'hbde598e1), .K8_C10_W4(32'hbdc176fd), .K8_C10_W5(32'hbd81a3a6), .K8_C10_W6(32'h3e1408df), .K8_C10_W7(32'hbd05b6a9), .K8_C10_W8(32'h3d7a7027), 
		.K8_C11_W0(32'h3da8134b), .K8_C11_W1(32'h3e09d78a), .K8_C11_W2(32'h3d280957), .K8_C11_W3(32'h3aef69d7), .K8_C11_W4(32'h3d1e9bf6), .K8_C11_W5(32'h3e05a629), .K8_C11_W6(32'h3c9282f5), .K8_C11_W7(32'h3d569456), .K8_C11_W8(32'hbe0151fd), 
		.K8_C12_W0(32'h3b8caffb), .K8_C12_W1(32'hbc955b8e), .K8_C12_W2(32'h3e168b40), .K8_C12_W3(32'h3d6d581c), .K8_C12_W4(32'h3df40868), .K8_C12_W5(32'hbde8ff83), .K8_C12_W6(32'h3de9a597), .K8_C12_W7(32'h3d4b81a3), .K8_C12_W8(32'hbdcdbe13), 
		.K8_C13_W0(32'h3dece77a), .K8_C13_W1(32'h3dc7c0da), .K8_C13_W2(32'h3d9f1260), .K8_C13_W3(32'h3e04eeff), .K8_C13_W4(32'h3da0c5ca), .K8_C13_W5(32'h3c4e35f3), .K8_C13_W6(32'h3d9b43c1), .K8_C13_W7(32'hbb50e551), .K8_C13_W8(32'hbdaa2544), 
		.K8_C14_W0(32'h3a757852), .K8_C14_W1(32'h3d05c049), .K8_C14_W2(32'hbd4cfe14), .K8_C14_W3(32'h3d7f63fc), .K8_C14_W4(32'hbd9c2aa2), .K8_C14_W5(32'hbd924906), .K8_C14_W6(32'h3daa3e28), .K8_C14_W7(32'hbd829e14), .K8_C14_W8(32'hbd66e293), 
		.K8_C15_W0(32'h3e0896ae), .K8_C15_W1(32'h3e0e4f16), .K8_C15_W2(32'h3d624544), .K8_C15_W3(32'hbe0e2265), .K8_C15_W4(32'h3db54f80), .K8_C15_W5(32'h3d0459db), .K8_C15_W6(32'hbd8dfb15), .K8_C15_W7(32'h3dece10a), .K8_C15_W8(32'hbd4449e3), 
		.K8_BIAS (32'h3cc37411),

		.K9_C0_W0(32'h3b15ca9b), .K9_C0_W1(32'hbd813b65), .K9_C0_W2(32'hbd43a9e6), .K9_C0_W3(32'h3d76ce7d), .K9_C0_W4(32'h3d804c65), .K9_C0_W5(32'hbdb73706), .K9_C0_W6(32'h3d0c6b2c), .K9_C0_W7(32'hbdc89c99), .K9_C0_W8(32'hbcb926f5), 
		.K9_C1_W0(32'h3db992be), .K9_C1_W1(32'h3d9caf13), .K9_C1_W2(32'hbdd2a4f6), .K9_C1_W3(32'hbd7622c6), .K9_C1_W4(32'hbd68c8ce), .K9_C1_W5(32'hbe05cf9d), .K9_C1_W6(32'hbe0533a7), .K9_C1_W7(32'h3ca12e80), .K9_C1_W8(32'h3d336035), 
		.K9_C2_W0(32'hbdfc475a), .K9_C2_W1(32'h3d56602c), .K9_C2_W2(32'h3e08e516), .K9_C2_W3(32'h3d4ddc81), .K9_C2_W4(32'h3d196b0f), .K9_C2_W5(32'hbe0ff03c), .K9_C2_W6(32'h3cee31b6), .K9_C2_W7(32'h3de44dd6), .K9_C2_W8(32'h3c6a200b), 
		.K9_C3_W0(32'hbdbce0d2), .K9_C3_W1(32'hbdc17885), .K9_C3_W2(32'hbccfd685), .K9_C3_W3(32'h3c94cf77), .K9_C3_W4(32'h3db5ae7a), .K9_C3_W5(32'h3d093d39), .K9_C3_W6(32'hbda68e64), .K9_C3_W7(32'hbe05cdb6), .K9_C3_W8(32'hbc9909cf), 
		.K9_C4_W0(32'hbc32d3a9), .K9_C4_W1(32'h3dc46f77), .K9_C4_W2(32'hbc8e5e1b), .K9_C4_W3(32'h3b3dd8e6), .K9_C4_W4(32'hbb363b30), .K9_C4_W5(32'hbd070808), .K9_C4_W6(32'h3da5597c), .K9_C4_W7(32'h3d33f8d5), .K9_C4_W8(32'hbc933a09), 
		.K9_C5_W0(32'h3dfd9ad2), .K9_C5_W1(32'hbe075fab), .K9_C5_W2(32'h3e18b318), .K9_C5_W3(32'h3ce5c083), .K9_C5_W4(32'h3be47d4e), .K9_C5_W5(32'h3ddc8312), .K9_C5_W6(32'hbd2c87ed), .K9_C5_W7(32'hbdc0cd5d), .K9_C5_W8(32'h3caf9f66), 
		.K9_C6_W0(32'hbcd6bc7d), .K9_C6_W1(32'h3c542ba2), .K9_C6_W2(32'h3c362ba2), .K9_C6_W3(32'hbcdeafde), .K9_C6_W4(32'hbddea7b4), .K9_C6_W5(32'h3cef55eb), .K9_C6_W6(32'h3ddf0e33), .K9_C6_W7(32'h3da2e708), .K9_C6_W8(32'h3db0b1f6), 
		.K9_C7_W0(32'h3de04ea8), .K9_C7_W1(32'hbd3f826c), .K9_C7_W2(32'hbddde051), .K9_C7_W3(32'h3e168900), .K9_C7_W4(32'h3d76fc3b), .K9_C7_W5(32'h3e0994e7), .K9_C7_W6(32'h3daeb8fe), .K9_C7_W7(32'h3dfcd91c), .K9_C7_W8(32'h3d86bf8a), 
		.K9_C8_W0(32'hbdf78afe), .K9_C8_W1(32'h3cd51e9f), .K9_C8_W2(32'hbe0c4d8c), .K9_C8_W3(32'hbd8ebe88), .K9_C8_W4(32'h3ddb2c38), .K9_C8_W5(32'h3e0c2bce), .K9_C8_W6(32'h3e0aec2c), .K9_C8_W7(32'hbd373e3e), .K9_C8_W8(32'hbcebe8b6), 
		.K9_C9_W0(32'h3dd5b749), .K9_C9_W1(32'h3d2a0457), .K9_C9_W2(32'h3d873f43), .K9_C9_W3(32'h3e13e787), .K9_C9_W4(32'h3df087dc), .K9_C9_W5(32'hbd908196), .K9_C9_W6(32'h3e1f7591), .K9_C9_W7(32'hbddfb2d5), .K9_C9_W8(32'h3e25956f), 
		.K9_C10_W0(32'h3e0c39ac), .K9_C10_W1(32'hbc8bd2d8), .K9_C10_W2(32'h3e004519), .K9_C10_W3(32'h3c591907), .K9_C10_W4(32'hbd8b7a6b), .K9_C10_W5(32'hbd841bcf), .K9_C10_W6(32'h3d732c83), .K9_C10_W7(32'hbcbfd89d), .K9_C10_W8(32'hbd720180), 
		.K9_C11_W0(32'hbe34ee8f), .K9_C11_W1(32'hbd36b270), .K9_C11_W2(32'hbde8b88a), .K9_C11_W3(32'hbde31e26), .K9_C11_W4(32'h3bdcc82b), .K9_C11_W5(32'hbd0bddb6), .K9_C11_W6(32'hbc9602e6), .K9_C11_W7(32'hbbefd07f), .K9_C11_W8(32'h3d4db713), 
		.K9_C12_W0(32'h3dd937d9), .K9_C12_W1(32'hbe1f870f), .K9_C12_W2(32'hbd29b09e), .K9_C12_W3(32'h3d5b06d5), .K9_C12_W4(32'hbcc78566), .K9_C12_W5(32'hbd2f79d7), .K9_C12_W6(32'h3bf0d43c), .K9_C12_W7(32'h3e0d1472), .K9_C12_W8(32'h3dc8bfe8), 
		.K9_C13_W0(32'hbdd995e5), .K9_C13_W1(32'h3dfc2b93), .K9_C13_W2(32'hbca4f4fa), .K9_C13_W3(32'h3d89a172), .K9_C13_W4(32'hbd51e682), .K9_C13_W5(32'h3c9ff5d2), .K9_C13_W6(32'hbd21697e), .K9_C13_W7(32'hbd8dfa93), .K9_C13_W8(32'hbdd9194f), 
		.K9_C14_W0(32'hbde59f61), .K9_C14_W1(32'h3e0ca896), .K9_C14_W2(32'h3debb508), .K9_C14_W3(32'h3d0fd85c), .K9_C14_W4(32'hbc579327), .K9_C14_W5(32'hbdef38d3), .K9_C14_W6(32'hbdf1e35f), .K9_C14_W7(32'hbcbc7e0c), .K9_C14_W8(32'hbde9f9de), 
		.K9_C15_W0(32'h3d2618b4), .K9_C15_W1(32'hbd2faa28), .K9_C15_W2(32'hbe215442), .K9_C15_W3(32'h3d8cd7b9), .K9_C15_W4(32'h3d191120), .K9_C15_W5(32'h3d3eb5fb), .K9_C15_W6(32'hbdb2301d), .K9_C15_W7(32'hbdfdb450), .K9_C15_W8(32'hbdb7c0aa), 
		.K9_BIAS (32'h3cd7bdbc),

		.K10_C0_W0(32'hbd135362), .K10_C0_W1(32'hbe070d6d), .K10_C0_W2(32'hbdad79eb), .K10_C0_W3(32'hbc39b5fc), .K10_C0_W4(32'hbc2ce1c1), .K10_C0_W5(32'h3dfb9cb0), .K10_C0_W6(32'h3ccea2e4), .K10_C0_W7(32'h3dea4393), .K10_C0_W8(32'h3dc1d2a5), 
		.K10_C1_W0(32'h3d17dc49), .K10_C1_W1(32'hbde843fc), .K10_C1_W2(32'hbcfe9ff3), .K10_C1_W3(32'h3dc50210), .K10_C1_W4(32'h3de4bf97), .K10_C1_W5(32'h3dbbc33a), .K10_C1_W6(32'hbd87a52d), .K10_C1_W7(32'hbda5760f), .K10_C1_W8(32'hbd44319c), 
		.K10_C2_W0(32'h3d993d33), .K10_C2_W1(32'hbdc6f3ab), .K10_C2_W2(32'h3dcd4cf0), .K10_C2_W3(32'hbd8559dd), .K10_C2_W4(32'h3e162dba), .K10_C2_W5(32'h3e31e6b1), .K10_C2_W6(32'hbdef8787), .K10_C2_W7(32'h3db0001a), .K10_C2_W8(32'hbd59ea0e), 
		.K10_C3_W0(32'h3d2b5b1d), .K10_C3_W1(32'hbddd0bd2), .K10_C3_W2(32'hbd278e49), .K10_C3_W3(32'hbcd077c7), .K10_C3_W4(32'hbda51886), .K10_C3_W5(32'h3d943e0a), .K10_C3_W6(32'hbe0b152b), .K10_C3_W7(32'h3dc3456c), .K10_C3_W8(32'hbd04c3be), 
		.K10_C4_W0(32'hbe2c8ce8), .K10_C4_W1(32'h3d364817), .K10_C4_W2(32'h3e02f205), .K10_C4_W3(32'hbc8a5538), .K10_C4_W4(32'hbd8f0193), .K10_C4_W5(32'hbdb9ae67), .K10_C4_W6(32'hbd8bbb47), .K10_C4_W7(32'h3d776f52), .K10_C4_W8(32'hbc27d60d), 
		.K10_C5_W0(32'hbd320761), .K10_C5_W1(32'h3debb0ae), .K10_C5_W2(32'hbdfe3217), .K10_C5_W3(32'h3d71e75e), .K10_C5_W4(32'hbdab1c7c), .K10_C5_W5(32'hbe21d25e), .K10_C5_W6(32'h3e03eeba), .K10_C5_W7(32'h3e1aec43), .K10_C5_W8(32'hbd375681), 
		.K10_C6_W0(32'hbe179606), .K10_C6_W1(32'hbc0156cd), .K10_C6_W2(32'hbdb2df02), .K10_C6_W3(32'hbdd119fd), .K10_C6_W4(32'hbd0bbc97), .K10_C6_W5(32'hbc01ae43), .K10_C6_W6(32'hbdf531bf), .K10_C6_W7(32'h3dad53e2), .K10_C6_W8(32'h3d9a3a03), 
		.K10_C7_W0(32'hbd56a811), .K10_C7_W1(32'hbdd132ca), .K10_C7_W2(32'hbe0f344a), .K10_C7_W3(32'hbd9f6b74), .K10_C7_W4(32'h3d953960), .K10_C7_W5(32'h3d6c405a), .K10_C7_W6(32'hbe098d96), .K10_C7_W7(32'h3b032578), .K10_C7_W8(32'h3d16fa2f), 
		.K10_C8_W0(32'hbd6751a9), .K10_C8_W1(32'h3d942108), .K10_C8_W2(32'h3d20206f), .K10_C8_W3(32'hbe07b589), .K10_C8_W4(32'hbdae354c), .K10_C8_W5(32'hbd036f0a), .K10_C8_W6(32'hbd707c28), .K10_C8_W7(32'hbda76a85), .K10_C8_W8(32'h3e2c05e7), 
		.K10_C9_W0(32'hbd39d13e), .K10_C9_W1(32'hbdf39326), .K10_C9_W2(32'hbd7d4f92), .K10_C9_W3(32'hba9fb95c), .K10_C9_W4(32'hbd4402ab), .K10_C9_W5(32'h3e15905f), .K10_C9_W6(32'hbd9068cb), .K10_C9_W7(32'hbc25db3a), .K10_C9_W8(32'h3e348fec), 
		.K10_C10_W0(32'hbceb5237), .K10_C10_W1(32'h3cfd9c1c), .K10_C10_W2(32'hbd9f8c4f), .K10_C10_W3(32'hbba7d794), .K10_C10_W4(32'h3d11b5d9), .K10_C10_W5(32'h3de258e1), .K10_C10_W6(32'h3dc7ae81), .K10_C10_W7(32'h3d90a867), .K10_C10_W8(32'hbe1d94a0), 
		.K10_C11_W0(32'h3d0e3932), .K10_C11_W1(32'hbdd85be2), .K10_C11_W2(32'hbd943c81), .K10_C11_W3(32'hbe09a8af), .K10_C11_W4(32'hb81b31f2), .K10_C11_W5(32'hbdb7bf2b), .K10_C11_W6(32'h3df3e45d), .K10_C11_W7(32'h3dbd30f4), .K10_C11_W8(32'hbd6fef1e), 
		.K10_C12_W0(32'hbdd2d27d), .K10_C12_W1(32'h3df569a4), .K10_C12_W2(32'hbcda86e0), .K10_C12_W3(32'hbd909695), .K10_C12_W4(32'hbe051a5b), .K10_C12_W5(32'hbe0a9d22), .K10_C12_W6(32'hbce08abc), .K10_C12_W7(32'hbe014f0d), .K10_C12_W8(32'hbd93577c), 
		.K10_C13_W0(32'hbc7bb7c3), .K10_C13_W1(32'hbe145707), .K10_C13_W2(32'h3dcc878f), .K10_C13_W3(32'hbc3669c4), .K10_C13_W4(32'h3d891474), .K10_C13_W5(32'hbdd2d7a4), .K10_C13_W6(32'h3d3c0ee6), .K10_C13_W7(32'hbd8791ba), .K10_C13_W8(32'h3d4a2f32), 
		.K10_C14_W0(32'hbd960cab), .K10_C14_W1(32'h3c0d83d2), .K10_C14_W2(32'hbdaaadeb), .K10_C14_W3(32'hbdb6e09b), .K10_C14_W4(32'hbdac3322), .K10_C14_W5(32'h3de8a803), .K10_C14_W6(32'h3d66503c), .K10_C14_W7(32'hbe1edc94), .K10_C14_W8(32'h3d861b2e), 
		.K10_C15_W0(32'h3a92cd42), .K10_C15_W1(32'hbd78b2c3), .K10_C15_W2(32'h3d3c119e), .K10_C15_W3(32'hbd46d7a1), .K10_C15_W4(32'hbc9bfe50), .K10_C15_W5(32'h3d7707f8), .K10_C15_W6(32'hbdda7d43), .K10_C15_W7(32'hbd93a011), .K10_C15_W8(32'h3da7b0b2), 
		.K10_BIAS (32'hbc87fe07),

		.K11_C0_W0(32'h3d38063a), .K11_C0_W1(32'hbccf5499), .K11_C0_W2(32'h3d93f450), .K11_C0_W3(32'hbe0ac36b), .K11_C0_W4(32'h3d718ef2), .K11_C0_W5(32'hbcd91902), .K11_C0_W6(32'hbd016f86), .K11_C0_W7(32'h3dd7713d), .K11_C0_W8(32'hbddabffc), 
		.K11_C1_W0(32'hbe197af1), .K11_C1_W1(32'hbdfc7a59), .K11_C1_W2(32'hbdd8829a), .K11_C1_W3(32'hbdbf47ad), .K11_C1_W4(32'h3905928e), .K11_C1_W5(32'h3def559e), .K11_C1_W6(32'hbc8565eb), .K11_C1_W7(32'h3c2c8bcb), .K11_C1_W8(32'hbd4c423c), 
		.K11_C2_W0(32'hbd7f9445), .K11_C2_W1(32'hbe0a3ec3), .K11_C2_W2(32'h3e008bbf), .K11_C2_W3(32'hbe175fc1), .K11_C2_W4(32'hbe041a23), .K11_C2_W5(32'h3d4d7852), .K11_C2_W6(32'hbd9b0c6f), .K11_C2_W7(32'hbd5d1a76), .K11_C2_W8(32'hbd91a05b), 
		.K11_C3_W0(32'h3e2c6441), .K11_C3_W1(32'hbdd6149b), .K11_C3_W2(32'hbda81f00), .K11_C3_W3(32'hbd2665ad), .K11_C3_W4(32'hbd70a6e9), .K11_C3_W5(32'hbc9fe5b9), .K11_C3_W6(32'h3e0d7417), .K11_C3_W7(32'h3e283bb4), .K11_C3_W8(32'h3d7105a7), 
		.K11_C4_W0(32'hbe430bb9), .K11_C4_W1(32'h3bdf09e4), .K11_C4_W2(32'h3d85c319), .K11_C4_W3(32'h3e121f4d), .K11_C4_W4(32'hbde6311e), .K11_C4_W5(32'hbd89bd2e), .K11_C4_W6(32'h3e06f346), .K11_C4_W7(32'h3dbc1dad), .K11_C4_W8(32'hbc6b8ec4), 
		.K11_C5_W0(32'hbdb991db), .K11_C5_W1(32'hbdca3d61), .K11_C5_W2(32'h3ddee1dc), .K11_C5_W3(32'hbdbf0407), .K11_C5_W4(32'hbcd76736), .K11_C5_W5(32'h3dc9aa78), .K11_C5_W6(32'hbd949ac5), .K11_C5_W7(32'h3d862f37), .K11_C5_W8(32'h3db2f00b), 
		.K11_C6_W0(32'hbba57122), .K11_C6_W1(32'hbd4c5e4c), .K11_C6_W2(32'hbd861017), .K11_C6_W3(32'h3d303f52), .K11_C6_W4(32'h3d9f97c1), .K11_C6_W5(32'hbceeee6e), .K11_C6_W6(32'hbd0c3640), .K11_C6_W7(32'h3dafe3c8), .K11_C6_W8(32'hbd765c28), 
		.K11_C7_W0(32'h3c245d63), .K11_C7_W1(32'h3cff6dea), .K11_C7_W2(32'hbd0824fe), .K11_C7_W3(32'h3e121bf6), .K11_C7_W4(32'h3d124154), .K11_C7_W5(32'hbdb83d38), .K11_C7_W6(32'hbc7cdafb), .K11_C7_W7(32'h3df2c1ef), .K11_C7_W8(32'hbdb425b4), 
		.K11_C8_W0(32'h3de14672), .K11_C8_W1(32'h3e0f3032), .K11_C8_W2(32'h3ca43352), .K11_C8_W3(32'h3d2bcbe2), .K11_C8_W4(32'h3d34267b), .K11_C8_W5(32'hbcd45192), .K11_C8_W6(32'h3ca89400), .K11_C8_W7(32'hbd08daee), .K11_C8_W8(32'hbd6af962), 
		.K11_C9_W0(32'hbe07c447), .K11_C9_W1(32'hbd3b90cc), .K11_C9_W2(32'hbd89047a), .K11_C9_W3(32'h3bce3179), .K11_C9_W4(32'h3c9b01b2), .K11_C9_W5(32'hbd564794), .K11_C9_W6(32'hbe0535fd), .K11_C9_W7(32'h3ddbea46), .K11_C9_W8(32'h3db0d627), 
		.K11_C10_W0(32'h3dde15fd), .K11_C10_W1(32'hbd402de5), .K11_C10_W2(32'h3d5f8e82), .K11_C10_W3(32'hbe12bdba), .K11_C10_W4(32'hbdb2f9dd), .K11_C10_W5(32'hbde8b23a), .K11_C10_W6(32'hbde0a1ee), .K11_C10_W7(32'h3db5342d), .K11_C10_W8(32'h3bdefca2), 
		.K11_C11_W0(32'h3d46ea5a), .K11_C11_W1(32'h3dd53985), .K11_C11_W2(32'hbde18358), .K11_C11_W3(32'h3dbe538c), .K11_C11_W4(32'hbce2e211), .K11_C11_W5(32'hbdfc9fc6), .K11_C11_W6(32'h3e01787c), .K11_C11_W7(32'h3da58140), .K11_C11_W8(32'hbda1945e), 
		.K11_C12_W0(32'h3dbd7255), .K11_C12_W1(32'hbd236842), .K11_C12_W2(32'h3e2036e8), .K11_C12_W3(32'hbdaa6014), .K11_C12_W4(32'hbc684582), .K11_C12_W5(32'h3da4ed5d), .K11_C12_W6(32'hbdbc4216), .K11_C12_W7(32'hbcb933dc), .K11_C12_W8(32'hbe205bb9), 
		.K11_C13_W0(32'h3d7bbbbd), .K11_C13_W1(32'h3d54e5bf), .K11_C13_W2(32'h3d9cf30a), .K11_C13_W3(32'hbdc07535), .K11_C13_W4(32'h3e08fc31), .K11_C13_W5(32'h3df7131c), .K11_C13_W6(32'h3d9db21f), .K11_C13_W7(32'hbe05af34), .K11_C13_W8(32'h3c24412e), 
		.K11_C14_W0(32'hbe0aaf49), .K11_C14_W1(32'hbddb64ca), .K11_C14_W2(32'h3d2c0570), .K11_C14_W3(32'h3c62f135), .K11_C14_W4(32'h3ddffd3d), .K11_C14_W5(32'h3dc89d97), .K11_C14_W6(32'h3b0d09bd), .K11_C14_W7(32'h3e41980b), .K11_C14_W8(32'hbda790ff), 
		.K11_C15_W0(32'hbdf93d49), .K11_C15_W1(32'h3dfbe7a2), .K11_C15_W2(32'h3dd21c85), .K11_C15_W3(32'hbe10da01), .K11_C15_W4(32'h3abc35cb), .K11_C15_W5(32'hbdce9a41), .K11_C15_W6(32'h3e1f548d), .K11_C15_W7(32'h3d9ea6cb), .K11_C15_W8(32'hbd87475d), 
		.K11_BIAS (32'hbd19e8c5),

		.K12_C0_W0(32'hbc1ff207), .K12_C0_W1(32'hbbe856ad), .K12_C0_W2(32'h3e130eaa), .K12_C0_W3(32'h3d1b75fe), .K12_C0_W4(32'hbe25d687), .K12_C0_W5(32'hbc9fc80b), .K12_C0_W6(32'hbdafb8e4), .K12_C0_W7(32'h3de7be7d), .K12_C0_W8(32'hbd049ab1), 
		.K12_C1_W0(32'h3b0d77ee), .K12_C1_W1(32'hbe0ef315), .K12_C1_W2(32'h3c0491c7), .K12_C1_W3(32'hbe23b548), .K12_C1_W4(32'hbdb6a948), .K12_C1_W5(32'h3d1e90fa), .K12_C1_W6(32'hbe2d5c89), .K12_C1_W7(32'h3deca442), .K12_C1_W8(32'h3d191903), 
		.K12_C2_W0(32'h3d739d7d), .K12_C2_W1(32'hbdbf0bca), .K12_C2_W2(32'hbd54a8b9), .K12_C2_W3(32'h3e1265d3), .K12_C2_W4(32'h3df31f22), .K12_C2_W5(32'hbce60da8), .K12_C2_W6(32'hbdccca74), .K12_C2_W7(32'hbbe4ef09), .K12_C2_W8(32'hbd848126), 
		.K12_C3_W0(32'h3d05b537), .K12_C3_W1(32'hbc886954), .K12_C3_W2(32'hbcceabac), .K12_C3_W3(32'h3db7bb8d), .K12_C3_W4(32'hbb56bd78), .K12_C3_W5(32'hbd3e91c8), .K12_C3_W6(32'hbc14605f), .K12_C3_W7(32'h3db1dba3), .K12_C3_W8(32'hbdb9565b), 
		.K12_C4_W0(32'hbdaf2358), .K12_C4_W1(32'h3d6b7c5a), .K12_C4_W2(32'h3d481307), .K12_C4_W3(32'hbe139ab6), .K12_C4_W4(32'hbe20a0e1), .K12_C4_W5(32'hbd041468), .K12_C4_W6(32'h3c4961f3), .K12_C4_W7(32'h3d0964f5), .K12_C4_W8(32'hbd7266fd), 
		.K12_C5_W0(32'hbcb91f63), .K12_C5_W1(32'hbc9e252f), .K12_C5_W2(32'hbe052955), .K12_C5_W3(32'h3db03e9e), .K12_C5_W4(32'h3b230945), .K12_C5_W5(32'h3d7b7a73), .K12_C5_W6(32'hbd91d414), .K12_C5_W7(32'hbdd7724f), .K12_C5_W8(32'hbb20defe), 
		.K12_C6_W0(32'h3be09de5), .K12_C6_W1(32'h3d25fc34), .K12_C6_W2(32'hbd46e625), .K12_C6_W3(32'h3e08e596), .K12_C6_W4(32'h3dd75b99), .K12_C6_W5(32'h3da0a658), .K12_C6_W6(32'h3c9ee05a), .K12_C6_W7(32'h3dd26745), .K12_C6_W8(32'hbd2023c7), 
		.K12_C7_W0(32'h3c9e73ab), .K12_C7_W1(32'hbd325600), .K12_C7_W2(32'h3de0d952), .K12_C7_W3(32'hbdaf7714), .K12_C7_W4(32'hbe0121d8), .K12_C7_W5(32'hbd4943a0), .K12_C7_W6(32'hbd44fe99), .K12_C7_W7(32'h3df78884), .K12_C7_W8(32'hbd0684c1), 
		.K12_C8_W0(32'h3c167d4d), .K12_C8_W1(32'h3be06741), .K12_C8_W2(32'hbda268d8), .K12_C8_W3(32'hbdc19685), .K12_C8_W4(32'h3e0f70d3), .K12_C8_W5(32'h3c574696), .K12_C8_W6(32'hbdaa3fdc), .K12_C8_W7(32'h3dafcce0), .K12_C8_W8(32'hbbe79f93), 
		.K12_C9_W0(32'hb929b794), .K12_C9_W1(32'hbdb95183), .K12_C9_W2(32'h3cd30499), .K12_C9_W3(32'h3dad4139), .K12_C9_W4(32'h3cec4906), .K12_C9_W5(32'hbdbe6ebe), .K12_C9_W6(32'h3d833c50), .K12_C9_W7(32'h3d6eb6d5), .K12_C9_W8(32'hbd072f88), 
		.K12_C10_W0(32'hbde4dc12), .K12_C10_W1(32'hbb03858d), .K12_C10_W2(32'hbe110cbf), .K12_C10_W3(32'h3d29e824), .K12_C10_W4(32'h3ca8a73e), .K12_C10_W5(32'h3c8c0d95), .K12_C10_W6(32'hbdea7061), .K12_C10_W7(32'hbd989069), .K12_C10_W8(32'h3dd29fb7), 
		.K12_C11_W0(32'h3ae89367), .K12_C11_W1(32'h3ccd93f4), .K12_C11_W2(32'h3d2b6b35), .K12_C11_W3(32'hbdf2f349), .K12_C11_W4(32'hbd81b240), .K12_C11_W5(32'hbe014aa6), .K12_C11_W6(32'hbb827c74), .K12_C11_W7(32'hbd6849f6), .K12_C11_W8(32'h3c22ad10), 
		.K12_C12_W0(32'h3da05dec), .K12_C12_W1(32'hbd635fd3), .K12_C12_W2(32'hbdf66f7f), .K12_C12_W3(32'h3e1185dd), .K12_C12_W4(32'h3d2b11a0), .K12_C12_W5(32'hbd71a48b), .K12_C12_W6(32'h3d850156), .K12_C12_W7(32'h3cff9fa6), .K12_C12_W8(32'hbcdd000c), 
		.K12_C13_W0(32'hbdefedd3), .K12_C13_W1(32'hbdcf5907), .K12_C13_W2(32'hbc90e147), .K12_C13_W3(32'hbde3d5fc), .K12_C13_W4(32'hbd7c5f6f), .K12_C13_W5(32'hbcdb9ae0), .K12_C13_W6(32'h3ca7020f), .K12_C13_W7(32'hbc9c063f), .K12_C13_W8(32'hbbcfab7c), 
		.K12_C14_W0(32'hbdad8bd3), .K12_C14_W1(32'h3d7c706b), .K12_C14_W2(32'h3d0793a3), .K12_C14_W3(32'hbd89a646), .K12_C14_W4(32'hbd944462), .K12_C14_W5(32'hbe10d3ee), .K12_C14_W6(32'hbc91eb70), .K12_C14_W7(32'hbdfa8b5c), .K12_C14_W8(32'hbdb03955), 
		.K12_C15_W0(32'h3d2f10c5), .K12_C15_W1(32'hbc9cdeaa), .K12_C15_W2(32'h3c6f47fe), .K12_C15_W3(32'hbd991625), .K12_C15_W4(32'hbd19f21b), .K12_C15_W5(32'hbcd789b1), .K12_C15_W6(32'h3deceae7), .K12_C15_W7(32'h3d79447c), .K12_C15_W8(32'hbdebe38e), 
		.K12_BIAS (32'hbd06c3fb),

		.K13_C0_W0(32'hbdcd89d0), .K13_C0_W1(32'h3c19c698), .K13_C0_W2(32'h3c209b09), .K13_C0_W3(32'hbcaee71f), .K13_C0_W4(32'h3d878b49), .K13_C0_W5(32'hbe301773), .K13_C0_W6(32'h3d78f3ad), .K13_C0_W7(32'hbe1c5f97), .K13_C0_W8(32'h3dd91378), 
		.K13_C1_W0(32'h3df42b66), .K13_C1_W1(32'h3db582ed), .K13_C1_W2(32'h3dab79f9), .K13_C1_W3(32'hbd3605b0), .K13_C1_W4(32'h3dafdf9a), .K13_C1_W5(32'hbe0d3b1a), .K13_C1_W6(32'h3de96857), .K13_C1_W7(32'hbe1e9309), .K13_C1_W8(32'hbd8bb712), 
		.K13_C2_W0(32'h3e0937ab), .K13_C2_W1(32'h3d0cd4e8), .K13_C2_W2(32'hbe1a5205), .K13_C2_W3(32'hbda88a07), .K13_C2_W4(32'h3c876d60), .K13_C2_W5(32'hbd2417e7), .K13_C2_W6(32'hbd716464), .K13_C2_W7(32'h3cc8f507), .K13_C2_W8(32'h3da404f9), 
		.K13_C3_W0(32'hbdb16eb7), .K13_C3_W1(32'h3daae282), .K13_C3_W2(32'hbe048164), .K13_C3_W3(32'h3e018dab), .K13_C3_W4(32'h3e0ef81e), .K13_C3_W5(32'h3e328300), .K13_C3_W6(32'h3de39a32), .K13_C3_W7(32'hbe11ec4d), .K13_C3_W8(32'h3d561ed1), 
		.K13_C4_W0(32'hbd7bb5e4), .K13_C4_W1(32'hbdb2b619), .K13_C4_W2(32'hbcb5954f), .K13_C4_W3(32'h3c85f83c), .K13_C4_W4(32'h3d148506), .K13_C4_W5(32'h3e02d29a), .K13_C4_W6(32'hbe05d87d), .K13_C4_W7(32'hbe21a246), .K13_C4_W8(32'h3b8aaa1c), 
		.K13_C5_W0(32'h3dd3aa4d), .K13_C5_W1(32'h3dba7341), .K13_C5_W2(32'h3e12c639), .K13_C5_W3(32'h3e58f340), .K13_C5_W4(32'h3dd5b106), .K13_C5_W5(32'hbd9c6f3b), .K13_C5_W6(32'hbd3d3d01), .K13_C5_W7(32'h3da89e57), .K13_C5_W8(32'h3ca3718f), 
		.K13_C6_W0(32'h3e011840), .K13_C6_W1(32'hbcbc31be), .K13_C6_W2(32'h3e118cc7), .K13_C6_W3(32'hbdb599b5), .K13_C6_W4(32'h3d663b97), .K13_C6_W5(32'h3cb51ef8), .K13_C6_W6(32'h3da07f97), .K13_C6_W7(32'h3d222ea6), .K13_C6_W8(32'h3e10c7fa), 
		.K13_C7_W0(32'h3e069efb), .K13_C7_W1(32'hbcd741d9), .K13_C7_W2(32'h3e0f5a57), .K13_C7_W3(32'hbcca4615), .K13_C7_W4(32'hbcd41f17), .K13_C7_W5(32'h3d9df998), .K13_C7_W6(32'hbbdd8a4d), .K13_C7_W7(32'hbd1bded5), .K13_C7_W8(32'h3d07f351), 
		.K13_C8_W0(32'hbe371eeb), .K13_C8_W1(32'h3de06ce9), .K13_C8_W2(32'h3d2eee41), .K13_C8_W3(32'hbe18f58f), .K13_C8_W4(32'h3d25c330), .K13_C8_W5(32'hbdb13342), .K13_C8_W6(32'hbde4ce66), .K13_C8_W7(32'hbdff9573), .K13_C8_W8(32'hbcad8f79), 
		.K13_C9_W0(32'h3d6018ec), .K13_C9_W1(32'h3ccff646), .K13_C9_W2(32'h3d9d3408), .K13_C9_W3(32'h3d0806d7), .K13_C9_W4(32'hbd964213), .K13_C9_W5(32'h3d9d5f75), .K13_C9_W6(32'h3e025ee3), .K13_C9_W7(32'h3dd4ae1e), .K13_C9_W8(32'hbc988aca), 
		.K13_C10_W0(32'h3e047a90), .K13_C10_W1(32'hbd7f43fb), .K13_C10_W2(32'h3d2674bf), .K13_C10_W3(32'h3de8ab5a), .K13_C10_W4(32'hbd8d1bad), .K13_C10_W5(32'hbc057f99), .K13_C10_W6(32'h3c34c737), .K13_C10_W7(32'hbd8affc0), .K13_C10_W8(32'hbc2bd272), 
		.K13_C11_W0(32'hbe10b6d8), .K13_C11_W1(32'hbd3b7a72), .K13_C11_W2(32'hbb92d02b), .K13_C11_W3(32'hbdad60af), .K13_C11_W4(32'h3dad91bf), .K13_C11_W5(32'hbc9ca2c3), .K13_C11_W6(32'h3b56a309), .K13_C11_W7(32'h3dd50626), .K13_C11_W8(32'hbe0c26a5), 
		.K13_C12_W0(32'h3b73ea57), .K13_C12_W1(32'hbca4c5a1), .K13_C12_W2(32'hbd276002), .K13_C12_W3(32'h3dc89feb), .K13_C12_W4(32'h3c1267bf), .K13_C12_W5(32'hbc9a83d7), .K13_C12_W6(32'h3d9b1fae), .K13_C12_W7(32'hbddfc22d), .K13_C12_W8(32'h3db0a1f7), 
		.K13_C13_W0(32'hbd55beb6), .K13_C13_W1(32'hbdcecfbd), .K13_C13_W2(32'h3d73cee0), .K13_C13_W3(32'hbc92b907), .K13_C13_W4(32'hbdd5fa5d), .K13_C13_W5(32'hbdffe64d), .K13_C13_W6(32'h3d2ac9e7), .K13_C13_W7(32'h3c89ed4e), .K13_C13_W8(32'h3d0e76ac), 
		.K13_C14_W0(32'h3de7416c), .K13_C14_W1(32'h3e0955ed), .K13_C14_W2(32'hbe05500f), .K13_C14_W3(32'h3d98bec2), .K13_C14_W4(32'hbd5f12e8), .K13_C14_W5(32'hbd6212f9), .K13_C14_W6(32'h3c4868d2), .K13_C14_W7(32'hbe049246), .K13_C14_W8(32'h3dfcc3b5), 
		.K13_C15_W0(32'hbdf6a16f), .K13_C15_W1(32'hbc50c831), .K13_C15_W2(32'h3da1bcf8), .K13_C15_W3(32'h3debc958), .K13_C15_W4(32'h3dbac864), .K13_C15_W5(32'hbde30d46), .K13_C15_W6(32'hbc23c0cf), .K13_C15_W7(32'hbe2a1378), .K13_C15_W8(32'h3df4b2ed), 
		.K13_BIAS (32'h3d5311c3),

		.K14_C0_W0(32'hbd4476a5), .K14_C0_W1(32'hbdbc3407), .K14_C0_W2(32'hbdb4e10a), .K14_C0_W3(32'h3e44ea3f), .K14_C0_W4(32'hbd66a974), .K14_C0_W5(32'h3e062bc5), .K14_C0_W6(32'h3e2d55c9), .K14_C0_W7(32'h3cc3a2f8), .K14_C0_W8(32'h3e3c4639), 
		.K14_C1_W0(32'hbe1c8233), .K14_C1_W1(32'h3d73e831), .K14_C1_W2(32'h3d743af2), .K14_C1_W3(32'hbd8bc6ea), .K14_C1_W4(32'h3d23a1ef), .K14_C1_W5(32'hbdd99457), .K14_C1_W6(32'h3d3efc61), .K14_C1_W7(32'hbd9bbc6b), .K14_C1_W8(32'hbd4267fc), 
		.K14_C2_W0(32'h3c3ab8dc), .K14_C2_W1(32'hbd0db947), .K14_C2_W2(32'h3d1b7567), .K14_C2_W3(32'hbe0dec88), .K14_C2_W4(32'h3ddb03b7), .K14_C2_W5(32'h3dd1f48f), .K14_C2_W6(32'hbd438b65), .K14_C2_W7(32'hbc52ca63), .K14_C2_W8(32'h3d3392d8), 
		.K14_C3_W0(32'hbd872e7c), .K14_C3_W1(32'hbda5756d), .K14_C3_W2(32'h3d4c5231), .K14_C3_W3(32'h3de3ac11), .K14_C3_W4(32'hbdefff64), .K14_C3_W5(32'h3ccb3fba), .K14_C3_W6(32'hbdf366d0), .K14_C3_W7(32'h3d59534a), .K14_C3_W8(32'hbddc29d4), 
		.K14_C4_W0(32'hbddf719b), .K14_C4_W1(32'hbd0a9967), .K14_C4_W2(32'h3d86b252), .K14_C4_W3(32'h3dfb853b), .K14_C4_W4(32'h3dd463d2), .K14_C4_W5(32'h3de1cc2b), .K14_C4_W6(32'hbb25b54a), .K14_C4_W7(32'hbbb18ab6), .K14_C4_W8(32'h3d153762), 
		.K14_C5_W0(32'h3c545113), .K14_C5_W1(32'h3d5dffd5), .K14_C5_W2(32'hba94b2f3), .K14_C5_W3(32'h3d7f72e8), .K14_C5_W4(32'h3d3da5ca), .K14_C5_W5(32'h3d8120b1), .K14_C5_W6(32'h3cc66be9), .K14_C5_W7(32'h3e002ce4), .K14_C5_W8(32'hbc231f31), 
		.K14_C6_W0(32'h3df38a40), .K14_C6_W1(32'h3c0ce6ec), .K14_C6_W2(32'hbdcf3e66), .K14_C6_W3(32'hbd8d0e82), .K14_C6_W4(32'h3c94f738), .K14_C6_W5(32'hbda668fd), .K14_C6_W6(32'hbd31586c), .K14_C6_W7(32'hbd86a40c), .K14_C6_W8(32'h3d58fc37), 
		.K14_C7_W0(32'h3bd53b0c), .K14_C7_W1(32'h3d0fc88d), .K14_C7_W2(32'hbafebf23), .K14_C7_W3(32'hbdc2bd5c), .K14_C7_W4(32'hbe16c116), .K14_C7_W5(32'hbdf3820c), .K14_C7_W6(32'hbd6ae2ac), .K14_C7_W7(32'h3dfdd02c), .K14_C7_W8(32'hbdf00d43), 
		.K14_C8_W0(32'h3d95341c), .K14_C8_W1(32'hbd89c900), .K14_C8_W2(32'h3c192b42), .K14_C8_W3(32'h3d57d5b2), .K14_C8_W4(32'h3d9208bc), .K14_C8_W5(32'hbd7fd522), .K14_C8_W6(32'h3db183fd), .K14_C8_W7(32'h3d903ea3), .K14_C8_W8(32'hbd00252d), 
		.K14_C9_W0(32'hbdb458fb), .K14_C9_W1(32'hbdcb0afe), .K14_C9_W2(32'h3c9d4414), .K14_C9_W3(32'h3da9f615), .K14_C9_W4(32'h3d5f6501), .K14_C9_W5(32'h3e01cbf1), .K14_C9_W6(32'h3d1b6c3b), .K14_C9_W7(32'hbd72d75d), .K14_C9_W8(32'hbe06c3ee), 
		.K14_C10_W0(32'hbd222a3a), .K14_C10_W1(32'hbe10a14e), .K14_C10_W2(32'h3d6e2b54), .K14_C10_W3(32'hbe34fd12), .K14_C10_W4(32'hbd8603b9), .K14_C10_W5(32'h3df66ef8), .K14_C10_W6(32'hbcf84e51), .K14_C10_W7(32'h3de45de8), .K14_C10_W8(32'h3dbf0d7d), 
		.K14_C11_W0(32'h3d0faaf2), .K14_C11_W1(32'h3e35a3af), .K14_C11_W2(32'hbd86fd78), .K14_C11_W3(32'hbcb1c432), .K14_C11_W4(32'hbe2a1382), .K14_C11_W5(32'hbe1cad7c), .K14_C11_W6(32'hbc94b3e8), .K14_C11_W7(32'h3d720a6e), .K14_C11_W8(32'hbdf15253), 
		.K14_C12_W0(32'hbdaf9951), .K14_C12_W1(32'h3d0c1c4f), .K14_C12_W2(32'hbdc9cfd4), .K14_C12_W3(32'hbd6d76e8), .K14_C12_W4(32'hbd533e4e), .K14_C12_W5(32'hbcf609a1), .K14_C12_W6(32'h3dd2b366), .K14_C12_W7(32'h3c9cb436), .K14_C12_W8(32'hbc96cc57), 
		.K14_C13_W0(32'h3e207dc5), .K14_C13_W1(32'h3d9d8b3a), .K14_C13_W2(32'h3ddf2711), .K14_C13_W3(32'hbd788f44), .K14_C13_W4(32'h3e2fcc7e), .K14_C13_W5(32'hbcd8cb42), .K14_C13_W6(32'hbd505389), .K14_C13_W7(32'hbcc46d99), .K14_C13_W8(32'hbd957a00), 
		.K14_C14_W0(32'hbd844706), .K14_C14_W1(32'hbde25460), .K14_C14_W2(32'hbd5c09d6), .K14_C14_W3(32'h3cf8a147), .K14_C14_W4(32'h3d8b2e17), .K14_C14_W5(32'hbd4d8b30), .K14_C14_W6(32'h3d92faa1), .K14_C14_W7(32'hbcb50820), .K14_C14_W8(32'h3ce02b21), 
		.K14_C15_W0(32'h3d6cb75e), .K14_C15_W1(32'hbd2e9eb6), .K14_C15_W2(32'hbe112920), .K14_C15_W3(32'h3d9cba8b), .K14_C15_W4(32'hbda8018b), .K14_C15_W5(32'hbdf4c193), .K14_C15_W6(32'hbc7c6e04), .K14_C15_W7(32'h3da311f7), .K14_C15_W8(32'h3de61999), 
		.K14_BIAS (32'hbcbfcc1a),

		.K15_C0_W0(32'h3cb6f2a5), .K15_C0_W1(32'h3da86ca2), .K15_C0_W2(32'h3d408298), .K15_C0_W3(32'h3cc70d23), .K15_C0_W4(32'h3d410b08), .K15_C0_W5(32'h3d28e676), .K15_C0_W6(32'hbd151632), .K15_C0_W7(32'h3dba7104), .K15_C0_W8(32'hbd9487ea), 
		.K15_C1_W0(32'h3ccb85d6), .K15_C1_W1(32'h3d9e9d1e), .K15_C1_W2(32'h3b90239b), .K15_C1_W3(32'h3d9e36e8), .K15_C1_W4(32'h3d8ba2b0), .K15_C1_W5(32'hbd860b4c), .K15_C1_W6(32'hbdfbb61e), .K15_C1_W7(32'hbd93c8f0), .K15_C1_W8(32'hbe0d3a12), 
		.K15_C2_W0(32'hbd8b3652), .K15_C2_W1(32'hbe093bad), .K15_C2_W2(32'hbe01bb33), .K15_C2_W3(32'h3d83e87e), .K15_C2_W4(32'h3dc6a7a0), .K15_C2_W5(32'hbd179be1), .K15_C2_W6(32'h3d92fa76), .K15_C2_W7(32'hbe178233), .K15_C2_W8(32'hbe130b89), 
		.K15_C3_W0(32'h3db2f4ae), .K15_C3_W1(32'h3cc54523), .K15_C3_W2(32'hbda8fb4f), .K15_C3_W3(32'h3e08b889), .K15_C3_W4(32'hbcd3c74d), .K15_C3_W5(32'hbe02879d), .K15_C3_W6(32'h3e18f24e), .K15_C3_W7(32'hbdc18665), .K15_C3_W8(32'hbdcabec5), 
		.K15_C4_W0(32'h3d0c9d56), .K15_C4_W1(32'h3b954f68), .K15_C4_W2(32'h3ce93364), .K15_C4_W3(32'h3c9954f1), .K15_C4_W4(32'h3ce8a720), .K15_C4_W5(32'h3d28166a), .K15_C4_W6(32'hbe02d0dc), .K15_C4_W7(32'h3d8a06c6), .K15_C4_W8(32'h3d23ac30), 
		.K15_C5_W0(32'hbdb51fcb), .K15_C5_W1(32'h3d2f7422), .K15_C5_W2(32'hbe0731c1), .K15_C5_W3(32'h3d38888d), .K15_C5_W4(32'h3db1ceff), .K15_C5_W5(32'h3de8cbdc), .K15_C5_W6(32'hbdab6d63), .K15_C5_W7(32'hbd7501b6), .K15_C5_W8(32'h3d886dd4), 
		.K15_C6_W0(32'h3d120d9e), .K15_C6_W1(32'hbc110f52), .K15_C6_W2(32'h3cf6e72e), .K15_C6_W3(32'h3dec7a5c), .K15_C6_W4(32'h3d552968), .K15_C6_W5(32'h3d9c1508), .K15_C6_W6(32'hbc68865e), .K15_C6_W7(32'h3dd5ae3c), .K15_C6_W8(32'h3b1de0b3), 
		.K15_C7_W0(32'h3a9b0d84), .K15_C7_W1(32'h3d390e2a), .K15_C7_W2(32'h3cbc9604), .K15_C7_W3(32'hbd539e95), .K15_C7_W4(32'hbc0255ad), .K15_C7_W5(32'h3d223b7f), .K15_C7_W6(32'h3e07578d), .K15_C7_W7(32'hbe1c5b44), .K15_C7_W8(32'h3c661fb3), 
		.K15_C8_W0(32'h3e1a6b3a), .K15_C8_W1(32'hbe114996), .K15_C8_W2(32'hbdd6292e), .K15_C8_W3(32'h3c87acc2), .K15_C8_W4(32'hbdfeddff), .K15_C8_W5(32'h3d2880a5), .K15_C8_W6(32'h3d1d8f8b), .K15_C8_W7(32'h3dbe9b3e), .K15_C8_W8(32'hbd138bad), 
		.K15_C9_W0(32'h3dc4a3ca), .K15_C9_W1(32'hbb782a62), .K15_C9_W2(32'hbda0701b), .K15_C9_W3(32'hbe0da076), .K15_C9_W4(32'h3c865d74), .K15_C9_W5(32'h3ce590d6), .K15_C9_W6(32'h3d390184), .K15_C9_W7(32'h3da6c088), .K15_C9_W8(32'h3e334aca), 
		.K15_C10_W0(32'hbb2c65f2), .K15_C10_W1(32'hbdbf6d97), .K15_C10_W2(32'h3d1b8669), .K15_C10_W3(32'hbe0289fb), .K15_C10_W4(32'h3daf628e), .K15_C10_W5(32'h3de70499), .K15_C10_W6(32'hbd7b47b6), .K15_C10_W7(32'h3dbca9cd), .K15_C10_W8(32'hbe0ad9b2), 
		.K15_C11_W0(32'h3dc29539), .K15_C11_W1(32'h3d407411), .K15_C11_W2(32'h3dd0cbf6), .K15_C11_W3(32'hbd199639), .K15_C11_W4(32'hbd25e239), .K15_C11_W5(32'hbcbbbd71), .K15_C11_W6(32'hbdb4265a), .K15_C11_W7(32'hbdb2cca6), .K15_C11_W8(32'h3d034f37), 
		.K15_C12_W0(32'hbdd4e9dd), .K15_C12_W1(32'h3db78dc2), .K15_C12_W2(32'h3e156ebe), .K15_C12_W3(32'hbdcabd84), .K15_C12_W4(32'hbd66e84c), .K15_C12_W5(32'h3e1438f0), .K15_C12_W6(32'h3deea340), .K15_C12_W7(32'h3e065a63), .K15_C12_W8(32'h3e0ad178), 
		.K15_C13_W0(32'h3e0c3d14), .K15_C13_W1(32'h3c26db72), .K15_C13_W2(32'hbdd460c6), .K15_C13_W3(32'h3d571f6b), .K15_C13_W4(32'h3d3723d4), .K15_C13_W5(32'h3d9dd514), .K15_C13_W6(32'h3de99cdc), .K15_C13_W7(32'h3d86805a), .K15_C13_W8(32'h3c132236), 
		.K15_C14_W0(32'hbe18e0b0), .K15_C14_W1(32'h3d90fda5), .K15_C14_W2(32'h3de955f9), .K15_C14_W3(32'h3cc7384d), .K15_C14_W4(32'h3cbc76b0), .K15_C14_W5(32'h3cb407d4), .K15_C14_W6(32'h3d9f0210), .K15_C14_W7(32'hbd92a02c), .K15_C14_W8(32'hbcd132fe), 
		.K15_C15_W0(32'h3df0126c), .K15_C15_W1(32'hbd852ec6), .K15_C15_W2(32'hbdbcde3f), .K15_C15_W3(32'hbbd3afc3), .K15_C15_W4(32'hbdb55703), .K15_C15_W5(32'hbd3ec546), .K15_C15_W6(32'h3d1d6241), .K15_C15_W7(32'h3ccc4ffe), .K15_C15_W8(32'h3e0d7b9e), 
		.K15_BIAS (32'hbd3f6096)
		)
		block4_conv2(
		.clk(clk),
		.resetn(resetn),
		.data_valid_in(conv_valid_out_4_1),
		.data_in_0(conv_out_4_1[0]),
		.data_in_1(conv_out_4_1[1]),
		.data_in_2(conv_out_4_1[2]),
		.data_in_3(conv_out_4_1[3]),
		.data_in_4(conv_out_4_1[4]),
		.data_in_5(conv_out_4_1[5]),
		.data_in_6(conv_out_4_1[6]),
		.data_in_7(conv_out_4_1[7]),
		.data_in_8(conv_out_4_1[8]),
		.data_in_9(conv_out_4_1[9]),
		.data_in_10(conv_out_4_1[10]),
		.data_in_11(conv_out_4_1[11]),
		.data_in_12(conv_out_4_1[12]),
		.data_in_13(conv_out_4_1[13]),
		.data_in_14(conv_out_4_1[14]),
		.data_in_15(conv_out_4_1[15]),
		.data_out_conv_0(conv_out_4_2[0]),
		.data_out_conv_1(conv_out_4_2[1]),
		.data_out_conv_2(conv_out_4_2[2]),
		.data_out_conv_3(conv_out_4_2[3]),
		.data_out_conv_4(conv_out_4_2[4]),
		.data_out_conv_5(conv_out_4_2[5]),
		.data_out_conv_6(conv_out_4_2[6]),
		.data_out_conv_7(conv_out_4_2[7]),
		.data_out_conv_8(conv_out_4_2[8]),
		.data_out_conv_9(conv_out_4_2[9]),
		.data_out_conv_10(conv_out_4_2[10]),
		.data_out_conv_11(conv_out_4_2[11]),
		.data_out_conv_12(conv_out_4_2[12]),
		.data_out_conv_13(conv_out_4_2[13]),
		.data_out_conv_14(conv_out_4_2[14]),
		.data_out_conv_15(conv_out_4_2[15]),
		.valid_out_pixel(conv_valid_out_4_2),
		.done(done_conv_4_2)
		);




	conv3d_16_kernel_16_channel_size_3 #(
		.DATA_WIDTH(32),.IMG_WIDTH(WIDTH),.IMG_HEIGHT(HEIGHT),
		.K0_C0_W0(32'hbdd94a6e), .K0_C0_W1(32'hbd4d4a9b), .K0_C0_W2(32'h3d930002), .K0_C0_W3(32'h3d958da6), .K0_C0_W4(32'hbced3357), .K0_C0_W5(32'h3de849d7), .K0_C0_W6(32'hbc919109), .K0_C0_W7(32'hbd358e00), .K0_C0_W8(32'h3e2a90c0), 
		.K0_C1_W0(32'h3c04e4eb), .K0_C1_W1(32'h3d03fb71), .K0_C1_W2(32'h3b2150a8), .K0_C1_W3(32'h3dd784be), .K0_C1_W4(32'h3e143d0e), .K0_C1_W5(32'h3df3e84c), .K0_C1_W6(32'h3d5240a1), .K0_C1_W7(32'h3cb7ca58), .K0_C1_W8(32'hbdfdcacb), 
		.K0_C2_W0(32'hbda526f2), .K0_C2_W1(32'h3d0114bc), .K0_C2_W2(32'hbb22a55b), .K0_C2_W3(32'hbdb51a02), .K0_C2_W4(32'h3daf4757), .K0_C2_W5(32'h3d03962c), .K0_C2_W6(32'hbe01290b), .K0_C2_W7(32'hbae29a18), .K0_C2_W8(32'hbd95edbf), 
		.K0_C3_W0(32'h3d42f886), .K0_C3_W1(32'hbc8280de), .K0_C3_W2(32'h3d8ecc3d), .K0_C3_W3(32'hbbe2786e), .K0_C3_W4(32'h3d92ed91), .K0_C3_W5(32'hbd4ba88b), .K0_C3_W6(32'hbdd89e26), .K0_C3_W7(32'hbd9fc999), .K0_C3_W8(32'h3d256cfc), 
		.K0_C4_W0(32'hbe19bfab), .K0_C4_W1(32'hbdccb794), .K0_C4_W2(32'h3d3e1aa0), .K0_C4_W3(32'h3d6a27b5), .K0_C4_W4(32'hbdcd3550), .K0_C4_W5(32'hbe161eb7), .K0_C4_W6(32'hbda7863b), .K0_C4_W7(32'h3df52a5a), .K0_C4_W8(32'hbe01ab30), 
		.K0_C5_W0(32'h3d962341), .K0_C5_W1(32'hbd0d1d29), .K0_C5_W2(32'hbe1f1ed4), .K0_C5_W3(32'h3dc7620b), .K0_C5_W4(32'h3dc80785), .K0_C5_W5(32'h3db5cd57), .K0_C5_W6(32'h3b63833a), .K0_C5_W7(32'hbdd52638), .K0_C5_W8(32'h3b9ef94c), 
		.K0_C6_W0(32'hbdfe2f5e), .K0_C6_W1(32'hbbe1852c), .K0_C6_W2(32'hbc787490), .K0_C6_W3(32'h3c470016), .K0_C6_W4(32'hbcde98f0), .K0_C6_W5(32'h3de77a84), .K0_C6_W6(32'h3c6137ae), .K0_C6_W7(32'hbde03815), .K0_C6_W8(32'h3d10025f), 
		.K0_C7_W0(32'hbdaf0247), .K0_C7_W1(32'h3d8238a6), .K0_C7_W2(32'hbd96332c), .K0_C7_W3(32'hbd93bbe7), .K0_C7_W4(32'hbc498505), .K0_C7_W5(32'hbd116102), .K0_C7_W6(32'hbd464ab8), .K0_C7_W7(32'hbc20fd8d), .K0_C7_W8(32'hbd179e67), 
		.K0_C8_W0(32'hbca24056), .K0_C8_W1(32'hbd7dd687), .K0_C8_W2(32'h3e146d68), .K0_C8_W3(32'hbd9698ad), .K0_C8_W4(32'hbcbe30a9), .K0_C8_W5(32'h3d31568b), .K0_C8_W6(32'h3cf8054f), .K0_C8_W7(32'h3cdbed45), .K0_C8_W8(32'h3cf91695), 
		.K0_C9_W0(32'hbe0b96bd), .K0_C9_W1(32'h3d4496cb), .K0_C9_W2(32'hbdddce16), .K0_C9_W3(32'h3e2a73a6), .K0_C9_W4(32'hbb85e0ec), .K0_C9_W5(32'h3df22a04), .K0_C9_W6(32'h3e1521df), .K0_C9_W7(32'hbd51ac5d), .K0_C9_W8(32'h3ddbc710), 
		.K0_C10_W0(32'h3de9442b), .K0_C10_W1(32'hbd517117), .K0_C10_W2(32'h3d7bfb69), .K0_C10_W3(32'h3d16f8ff), .K0_C10_W4(32'hbe0a6b62), .K0_C10_W5(32'hbe13bf8f), .K0_C10_W6(32'hbdca0a51), .K0_C10_W7(32'h3ddc6061), .K0_C10_W8(32'h3cbab08e), 
		.K0_C11_W0(32'h3c2e4499), .K0_C11_W1(32'h3d3a439e), .K0_C11_W2(32'hbd3e2017), .K0_C11_W3(32'h3cf9ca0e), .K0_C11_W4(32'h3cc361f8), .K0_C11_W5(32'hba3f97e9), .K0_C11_W6(32'h3c70a499), .K0_C11_W7(32'hbdd98897), .K0_C11_W8(32'hbde8a2cf), 
		.K0_C12_W0(32'hbdabd44f), .K0_C12_W1(32'hbe1832be), .K0_C12_W2(32'hbd757ffe), .K0_C12_W3(32'hbdb530a8), .K0_C12_W4(32'h3c0ccd92), .K0_C12_W5(32'hbddd947d), .K0_C12_W6(32'h3c27ff3c), .K0_C12_W7(32'h3ccd3f04), .K0_C12_W8(32'hbc844491), 
		.K0_C13_W0(32'h3d1cb6cb), .K0_C13_W1(32'hbdc70f19), .K0_C13_W2(32'hbcb6976a), .K0_C13_W3(32'h3e128591), .K0_C13_W4(32'hbd422a22), .K0_C13_W5(32'hbdb85d37), .K0_C13_W6(32'h3e2c0338), .K0_C13_W7(32'h3d8bcde3), .K0_C13_W8(32'hbd9937b4), 
		.K0_C14_W0(32'hbd874e0f), .K0_C14_W1(32'hbe13fdf3), .K0_C14_W2(32'hbd5253c2), .K0_C14_W3(32'hbdf82150), .K0_C14_W4(32'hbd5b45a4), .K0_C14_W5(32'hbe1b7278), .K0_C14_W6(32'h3c08bd13), .K0_C14_W7(32'hbe00594c), .K0_C14_W8(32'hbe05c54c), 
		.K0_C15_W0(32'hbd7282e6), .K0_C15_W1(32'h3d24c317), .K0_C15_W2(32'hbd0d4429), .K0_C15_W3(32'h3dfbf347), .K0_C15_W4(32'h3cbe1835), .K0_C15_W5(32'hbde782dd), .K0_C15_W6(32'h3dcd4e5c), .K0_C15_W7(32'hbe064cf8), .K0_C15_W8(32'h3df43b8d), 
		.K0_BIAS (32'h3d1f9130),

		.K1_C0_W0(32'hbc3f913a), .K1_C0_W1(32'hbcca3705), .K1_C0_W2(32'hbcc712ad), .K1_C0_W3(32'hbd3892b9), .K1_C0_W4(32'h3b16dc3a), .K1_C0_W5(32'h3d39a07d), .K1_C0_W6(32'hbda38bd8), .K1_C0_W7(32'hbdd7b778), .K1_C0_W8(32'h3dbf4e2f), 
		.K1_C1_W0(32'h3e0abffa), .K1_C1_W1(32'h3b72ebc2), .K1_C1_W2(32'h3dfea044), .K1_C1_W3(32'h3e18ff72), .K1_C1_W4(32'hbd8ed635), .K1_C1_W5(32'h3db6c59d), .K1_C1_W6(32'h3e07538f), .K1_C1_W7(32'hbcbfd6de), .K1_C1_W8(32'hbd98258d), 
		.K1_C2_W0(32'h3deface8), .K1_C2_W1(32'hbb95500e), .K1_C2_W2(32'h3d6f00f9), .K1_C2_W3(32'h3dfa25d5), .K1_C2_W4(32'h3d8206db), .K1_C2_W5(32'hbd29c32f), .K1_C2_W6(32'h3e0e13ec), .K1_C2_W7(32'hbd759811), .K1_C2_W8(32'h3bcd871d), 
		.K1_C3_W0(32'hbda47039), .K1_C3_W1(32'hbcaa1e87), .K1_C3_W2(32'h3d2c4ab9), .K1_C3_W3(32'hbddb1857), .K1_C3_W4(32'hbd427db1), .K1_C3_W5(32'h3d9c34bc), .K1_C3_W6(32'hbe28384c), .K1_C3_W7(32'h3dbd06c3), .K1_C3_W8(32'hbd88d465), 
		.K1_C4_W0(32'h3d7dcd03), .K1_C4_W1(32'hbda16106), .K1_C4_W2(32'h3c11b698), .K1_C4_W3(32'h3cb9a376), .K1_C4_W4(32'hbd8aeafd), .K1_C4_W5(32'hbd84e1ba), .K1_C4_W6(32'h3e1779ee), .K1_C4_W7(32'hbd9d6947), .K1_C4_W8(32'h3e2a70f9), 
		.K1_C5_W0(32'h3e137a1d), .K1_C5_W1(32'hbdb6aae1), .K1_C5_W2(32'h3cbd752d), .K1_C5_W3(32'hbca286a0), .K1_C5_W4(32'h3d46fcf3), .K1_C5_W5(32'h3e3a93a2), .K1_C5_W6(32'hbd7bdd8d), .K1_C5_W7(32'h3d43c0e2), .K1_C5_W8(32'h3deb3084), 
		.K1_C6_W0(32'hbd97aeed), .K1_C6_W1(32'h3d38ad1f), .K1_C6_W2(32'h3da57d02), .K1_C6_W3(32'hbe17d6df), .K1_C6_W4(32'hbd9c50ab), .K1_C6_W5(32'h3d9fad5b), .K1_C6_W6(32'h3c3c983f), .K1_C6_W7(32'hbdbdba67), .K1_C6_W8(32'h3d0eabe4), 
		.K1_C7_W0(32'h3d92cc94), .K1_C7_W1(32'h3dcac556), .K1_C7_W2(32'hbdb34058), .K1_C7_W3(32'h3df01627), .K1_C7_W4(32'h3e22fb75), .K1_C7_W5(32'h3dbb4d13), .K1_C7_W6(32'h3dabd6bf), .K1_C7_W7(32'h3d84cfe6), .K1_C7_W8(32'h3ced07d0), 
		.K1_C8_W0(32'h3dd7da32), .K1_C8_W1(32'hbd59648b), .K1_C8_W2(32'h3d987477), .K1_C8_W3(32'hbd23e822), .K1_C8_W4(32'hbd2d52c7), .K1_C8_W5(32'hbe335a2e), .K1_C8_W6(32'hbdf7bf7a), .K1_C8_W7(32'hbe20d055), .K1_C8_W8(32'hbdc267d7), 
		.K1_C9_W0(32'hbbbdcd2d), .K1_C9_W1(32'hbce3af9c), .K1_C9_W2(32'hbd7e05ad), .K1_C9_W3(32'hbd1e53d0), .K1_C9_W4(32'h3d07cb8f), .K1_C9_W5(32'h3dffb331), .K1_C9_W6(32'h3df84410), .K1_C9_W7(32'h3dc07aa8), .K1_C9_W8(32'h3df12279), 
		.K1_C10_W0(32'h3df354ee), .K1_C10_W1(32'h3b8e1f26), .K1_C10_W2(32'h3c5c9f53), .K1_C10_W3(32'h3e123eed), .K1_C10_W4(32'h3db431b1), .K1_C10_W5(32'h3db83640), .K1_C10_W6(32'hbd2b4d0e), .K1_C10_W7(32'hbdda4363), .K1_C10_W8(32'h3d1849c1), 
		.K1_C11_W0(32'h3d36b824), .K1_C11_W1(32'h3d74e314), .K1_C11_W2(32'h3de2496c), .K1_C11_W3(32'hbccb11ff), .K1_C11_W4(32'h3d047372), .K1_C11_W5(32'hbd34bafd), .K1_C11_W6(32'h3cca62e4), .K1_C11_W7(32'h3dd0e7ac), .K1_C11_W8(32'hbd9f7fa4), 
		.K1_C12_W0(32'h3de2b42a), .K1_C12_W1(32'hbcd721bd), .K1_C12_W2(32'hbd80ac5f), .K1_C12_W3(32'hbd486835), .K1_C12_W4(32'hbca2338e), .K1_C12_W5(32'h3c469e40), .K1_C12_W6(32'h3d80c62b), .K1_C12_W7(32'h3d9ec17c), .K1_C12_W8(32'h3e12356b), 
		.K1_C13_W0(32'h3b8d8d4e), .K1_C13_W1(32'h3e1c0981), .K1_C13_W2(32'hbde285b1), .K1_C13_W3(32'h3d199aaa), .K1_C13_W4(32'h3e082d09), .K1_C13_W5(32'hbdc19adc), .K1_C13_W6(32'hbbb0203a), .K1_C13_W7(32'hbd662189), .K1_C13_W8(32'h3e222440), 
		.K1_C14_W0(32'h3da8ecf5), .K1_C14_W1(32'hbda360ab), .K1_C14_W2(32'h3d6be8a0), .K1_C14_W3(32'hbd297335), .K1_C14_W4(32'hbe0f54ef), .K1_C14_W5(32'h3d3786f7), .K1_C14_W6(32'h3e1837df), .K1_C14_W7(32'h3d8ca7de), .K1_C14_W8(32'hbd68054c), 
		.K1_C15_W0(32'h3dd174aa), .K1_C15_W1(32'h3d9e66c2), .K1_C15_W2(32'h3cdcce44), .K1_C15_W3(32'hbde5ea63), .K1_C15_W4(32'h3cebd381), .K1_C15_W5(32'hbdb75166), .K1_C15_W6(32'h3d0aa3e4), .K1_C15_W7(32'hbd96be96), .K1_C15_W8(32'hbd7355b9), 
		.K1_BIAS (32'h3c0a67a0),

		.K2_C0_W0(32'hbde2fb3e), .K2_C0_W1(32'h3dbc88d3), .K2_C0_W2(32'hbb922b77), .K2_C0_W3(32'h3e08be83), .K2_C0_W4(32'hbd941b29), .K2_C0_W5(32'h3d9e2083), .K2_C0_W6(32'h3cfa5894), .K2_C0_W7(32'h3c99c004), .K2_C0_W8(32'hbe01fc9e), 
		.K2_C1_W0(32'hbd925013), .K2_C1_W1(32'h3d2c4e31), .K2_C1_W2(32'h3c28d260), .K2_C1_W3(32'h3e1274ca), .K2_C1_W4(32'hbd86afdb), .K2_C1_W5(32'hbddcb834), .K2_C1_W6(32'h3d430935), .K2_C1_W7(32'hbc1a170f), .K2_C1_W8(32'hbbc372f1), 
		.K2_C2_W0(32'h3dc8df01), .K2_C2_W1(32'hbdb839ae), .K2_C2_W2(32'hbd9b4400), .K2_C2_W3(32'h3dea9bed), .K2_C2_W4(32'hbd13bb3a), .K2_C2_W5(32'hbd865802), .K2_C2_W6(32'h3d44ab2f), .K2_C2_W7(32'hbb9cb1f9), .K2_C2_W8(32'hbd53f2b1), 
		.K2_C3_W0(32'h3dc61274), .K2_C3_W1(32'h3c27e5c6), .K2_C3_W2(32'hbd9e7983), .K2_C3_W3(32'hbda07718), .K2_C3_W4(32'hbd7d4709), .K2_C3_W5(32'h3dc09d32), .K2_C3_W6(32'hbb4eb929), .K2_C3_W7(32'hbd2114bb), .K2_C3_W8(32'hbd99b3b7), 
		.K2_C4_W0(32'hbda9e036), .K2_C4_W1(32'h3d22196a), .K2_C4_W2(32'hbd56cf1c), .K2_C4_W3(32'hbc832cf3), .K2_C4_W4(32'h3d6764ab), .K2_C4_W5(32'h3e05af06), .K2_C4_W6(32'h3db81730), .K2_C4_W7(32'hbcdcf5ff), .K2_C4_W8(32'h3cfa7231), 
		.K2_C5_W0(32'h3ddffc82), .K2_C5_W1(32'hbdcc1756), .K2_C5_W2(32'hbdcf564b), .K2_C5_W3(32'h3d15efb2), .K2_C5_W4(32'hbda2890f), .K2_C5_W5(32'h3d854b61), .K2_C5_W6(32'hbb86a3b2), .K2_C5_W7(32'hbddf7771), .K2_C5_W8(32'hbd397cfd), 
		.K2_C6_W0(32'hbdb16fb5), .K2_C6_W1(32'h3c77be9b), .K2_C6_W2(32'h3dbe88f7), .K2_C6_W3(32'hbcee14ea), .K2_C6_W4(32'hbdcf3989), .K2_C6_W5(32'h3dfee5eb), .K2_C6_W6(32'hbd71b3d3), .K2_C6_W7(32'hbdb120c8), .K2_C6_W8(32'h3e0e393f), 
		.K2_C7_W0(32'h3c3ccc52), .K2_C7_W1(32'hbde5e489), .K2_C7_W2(32'hbdff11ee), .K2_C7_W3(32'hbd7909ce), .K2_C7_W4(32'hbded2c17), .K2_C7_W5(32'hbda559c3), .K2_C7_W6(32'hbe06a236), .K2_C7_W7(32'h3dec0356), .K2_C7_W8(32'h3d36fcf7), 
		.K2_C8_W0(32'h3d6e70ee), .K2_C8_W1(32'hbce4e2aa), .K2_C8_W2(32'hbd393732), .K2_C8_W3(32'h3da14cdd), .K2_C8_W4(32'h3d11558d), .K2_C8_W5(32'hbd1de2e6), .K2_C8_W6(32'h3e0fe63a), .K2_C8_W7(32'h3d5be307), .K2_C8_W8(32'hbdafff25), 
		.K2_C9_W0(32'hbd83e30b), .K2_C9_W1(32'h3ce18d51), .K2_C9_W2(32'hbd66d619), .K2_C9_W3(32'hbe1e9477), .K2_C9_W4(32'h3de17a5e), .K2_C9_W5(32'hbddb19c1), .K2_C9_W6(32'hbe212afc), .K2_C9_W7(32'hbcf97a08), .K2_C9_W8(32'h3db65834), 
		.K2_C10_W0(32'h3d42f26a), .K2_C10_W1(32'h3db03d56), .K2_C10_W2(32'hbd5d1b4a), .K2_C10_W3(32'h3dadb8e9), .K2_C10_W4(32'hbaa1f81b), .K2_C10_W5(32'h3e108de8), .K2_C10_W6(32'h3d71cb37), .K2_C10_W7(32'hbd5195fc), .K2_C10_W8(32'hbdf65716), 
		.K2_C11_W0(32'hbdd2c613), .K2_C11_W1(32'h3dddfadf), .K2_C11_W2(32'h3dd741fb), .K2_C11_W3(32'hbd3bc815), .K2_C11_W4(32'h3d2f4272), .K2_C11_W5(32'h3e04cd44), .K2_C11_W6(32'hbd8eab33), .K2_C11_W7(32'h3d8e325a), .K2_C11_W8(32'h3cc866f4), 
		.K2_C12_W0(32'h3cbcfe9f), .K2_C12_W1(32'hbd8b62d6), .K2_C12_W2(32'hbdcb7009), .K2_C12_W3(32'h3e009f34), .K2_C12_W4(32'hbd89cd7a), .K2_C12_W5(32'hbd8761ca), .K2_C12_W6(32'hbd25926b), .K2_C12_W7(32'h3dbec5b7), .K2_C12_W8(32'hbdc0145a), 
		.K2_C13_W0(32'h3e0c05fc), .K2_C13_W1(32'hbdb71401), .K2_C13_W2(32'h3dbfbbe8), .K2_C13_W3(32'h3db6b206), .K2_C13_W4(32'hbd336965), .K2_C13_W5(32'hbd4b4d89), .K2_C13_W6(32'hbe2603d0), .K2_C13_W7(32'hbe23a19a), .K2_C13_W8(32'hbae3400b), 
		.K2_C14_W0(32'hbd81c29e), .K2_C14_W1(32'h3c88ea94), .K2_C14_W2(32'h3de23cd9), .K2_C14_W3(32'hbdceec2a), .K2_C14_W4(32'hbdd087ca), .K2_C14_W5(32'h3d07f61a), .K2_C14_W6(32'h3de289ae), .K2_C14_W7(32'h3d105b84), .K2_C14_W8(32'h3e1ad24f), 
		.K2_C15_W0(32'hbe1ab88c), .K2_C15_W1(32'h3db9eac3), .K2_C15_W2(32'h3ccb8228), .K2_C15_W3(32'hbd90b9fe), .K2_C15_W4(32'hbda9a52e), .K2_C15_W5(32'h3ce56994), .K2_C15_W6(32'hbdac3d6a), .K2_C15_W7(32'hbd7a3d32), .K2_C15_W8(32'h3df534b6), 
		.K2_BIAS (32'h3bb6f9be),

		.K3_C0_W0(32'hbdb1a845), .K3_C0_W1(32'hbc882034), .K3_C0_W2(32'h3dd7caee), .K3_C0_W3(32'hbca230af), .K3_C0_W4(32'h3e19c5e1), .K3_C0_W5(32'h3e09c2f8), .K3_C0_W6(32'h3e30e805), .K3_C0_W7(32'h3e1062c6), .K3_C0_W8(32'h3d77def7), 
		.K3_C1_W0(32'h3cae7df8), .K3_C1_W1(32'h3bd9e45f), .K3_C1_W2(32'h3cc77926), .K3_C1_W3(32'h3d590c6d), .K3_C1_W4(32'hbd132969), .K3_C1_W5(32'hba87cc56), .K3_C1_W6(32'hbdf3b77c), .K3_C1_W7(32'h3d652564), .K3_C1_W8(32'h3decc70c), 
		.K3_C2_W0(32'hbe14811b), .K3_C2_W1(32'h3dd12c88), .K3_C2_W2(32'hbdd56108), .K3_C2_W3(32'hbdf06532), .K3_C2_W4(32'hbd44816b), .K3_C2_W5(32'h3db71dac), .K3_C2_W6(32'hbdf8f1f7), .K3_C2_W7(32'hbc8c11a6), .K3_C2_W8(32'hbda7bbc2), 
		.K3_C3_W0(32'h3dc7236c), .K3_C3_W1(32'hbca678c1), .K3_C3_W2(32'h3e03fb8a), .K3_C3_W3(32'hbdf3a795), .K3_C3_W4(32'h3b4c3505), .K3_C3_W5(32'hbd0bc072), .K3_C3_W6(32'h3c510a28), .K3_C3_W7(32'h3d3016c1), .K3_C3_W8(32'h3d016188), 
		.K3_C4_W0(32'hbd5f9afe), .K3_C4_W1(32'h3d88625b), .K3_C4_W2(32'h3dbc4702), .K3_C4_W3(32'h3dcdd31f), .K3_C4_W4(32'h3d809ce2), .K3_C4_W5(32'hbd33616d), .K3_C4_W6(32'h3cfc9aec), .K3_C4_W7(32'h3e148018), .K3_C4_W8(32'h3df032c6), 
		.K3_C5_W0(32'hbd96e114), .K3_C5_W1(32'h3d54b92e), .K3_C5_W2(32'hbd890eb3), .K3_C5_W3(32'h3dd696d0), .K3_C5_W4(32'hbdbe98d4), .K3_C5_W5(32'hbe1031bf), .K3_C5_W6(32'hbd2b2d35), .K3_C5_W7(32'hbd894a89), .K3_C5_W8(32'hbcbdaa55), 
		.K3_C6_W0(32'h3e0a9f28), .K3_C6_W1(32'h3e0a1a05), .K3_C6_W2(32'hbd301d17), .K3_C6_W3(32'hbe3a3ba7), .K3_C6_W4(32'hbd326af8), .K3_C6_W5(32'h3c3f5dcc), .K3_C6_W6(32'hbde744dc), .K3_C6_W7(32'h3d5dd969), .K3_C6_W8(32'hbe06261c), 
		.K3_C7_W0(32'hbd397409), .K3_C7_W1(32'hbce17b64), .K3_C7_W2(32'h3cc593c7), .K3_C7_W3(32'hbc8ec8c1), .K3_C7_W4(32'h3dccd4e1), .K3_C7_W5(32'h3d880669), .K3_C7_W6(32'hbd3aaad4), .K3_C7_W7(32'h3c3bfd24), .K3_C7_W8(32'h3d328ddd), 
		.K3_C8_W0(32'hbe110f3e), .K3_C8_W1(32'hbbacd4c1), .K3_C8_W2(32'hbcd67162), .K3_C8_W3(32'hbd2bae04), .K3_C8_W4(32'hbb8f3617), .K3_C8_W5(32'h3de2f4fc), .K3_C8_W6(32'hbdba19ef), .K3_C8_W7(32'hbd1e37d7), .K3_C8_W8(32'hbdd2d2e0), 
		.K3_C9_W0(32'h3c8b505d), .K3_C9_W1(32'h3dfb678a), .K3_C9_W2(32'h3c5b9a2c), .K3_C9_W3(32'hbde92ac4), .K3_C9_W4(32'hbe07dde8), .K3_C9_W5(32'hbca54ae6), .K3_C9_W6(32'hbd3de232), .K3_C9_W7(32'hbdb4276f), .K3_C9_W8(32'h3dec841b), 
		.K3_C10_W0(32'hbde443fd), .K3_C10_W1(32'hbdfea480), .K3_C10_W2(32'h3dd9d3be), .K3_C10_W3(32'h3d326b45), .K3_C10_W4(32'h3d31f52b), .K3_C10_W5(32'h3db11f09), .K3_C10_W6(32'h3c56e2e5), .K3_C10_W7(32'hbd4ca9f6), .K3_C10_W8(32'hbd07c4e4), 
		.K3_C11_W0(32'hbe0e5a1f), .K3_C11_W1(32'h3d6a9c5b), .K3_C11_W2(32'hbdf88461), .K3_C11_W3(32'h3df2ecc6), .K3_C11_W4(32'hbcce8a29), .K3_C11_W5(32'hbbd5e344), .K3_C11_W6(32'h3d509c1f), .K3_C11_W7(32'h3ad0445c), .K3_C11_W8(32'h3c6f6db4), 
		.K3_C12_W0(32'h3d792692), .K3_C12_W1(32'hbbd66923), .K3_C12_W2(32'h3dc7c733), .K3_C12_W3(32'h3c49db85), .K3_C12_W4(32'hbe11cc45), .K3_C12_W5(32'h3cd87f51), .K3_C12_W6(32'h3d42a07c), .K3_C12_W7(32'h3d3c87a0), .K3_C12_W8(32'hbda4a69e), 
		.K3_C13_W0(32'hbbc334e7), .K3_C13_W1(32'hbdf16c1d), .K3_C13_W2(32'h3dec4ca6), .K3_C13_W3(32'h3e411b97), .K3_C13_W4(32'hbd2e65c6), .K3_C13_W5(32'h3b8bd7f5), .K3_C13_W6(32'h3ddb63f3), .K3_C13_W7(32'h3db2f475), .K3_C13_W8(32'h3e11d7d5), 
		.K3_C14_W0(32'h3df25f52), .K3_C14_W1(32'h3de27d0e), .K3_C14_W2(32'h3ca42a45), .K3_C14_W3(32'hbdb7211f), .K3_C14_W4(32'hbdfaf661), .K3_C14_W5(32'h3e0756ca), .K3_C14_W6(32'h3e1b1c25), .K3_C14_W7(32'hbc0ff0e3), .K3_C14_W8(32'hbdc82a4e), 
		.K3_C15_W0(32'hbe4dcd34), .K3_C15_W1(32'hbdbcdda6), .K3_C15_W2(32'hbccabda9), .K3_C15_W3(32'hbcac0874), .K3_C15_W4(32'hbe11face), .K3_C15_W5(32'h3c126d48), .K3_C15_W6(32'hbd499e27), .K3_C15_W7(32'h3d4211af), .K3_C15_W8(32'hbe0ee97d), 
		.K3_BIAS (32'h3cf1e7bb),

		.K4_C0_W0(32'h3ce7e593), .K4_C0_W1(32'hbd6c5e85), .K4_C0_W2(32'hbd9dc2cb), .K4_C0_W3(32'h3ddfa7e9), .K4_C0_W4(32'h3de04746), .K4_C0_W5(32'hbd33a9f0), .K4_C0_W6(32'h3d0436b7), .K4_C0_W7(32'hbdc3e17a), .K4_C0_W8(32'h3d2d3f8b), 
		.K4_C1_W0(32'hbdc1fd6d), .K4_C1_W1(32'hbda82a38), .K4_C1_W2(32'h3afa5dde), .K4_C1_W3(32'h3c3516b0), .K4_C1_W4(32'hbd0d93fa), .K4_C1_W5(32'hbe0faab4), .K4_C1_W6(32'h3dae99b9), .K4_C1_W7(32'hbc28f0fb), .K4_C1_W8(32'hbda62a65), 
		.K4_C2_W0(32'hbd14b6d3), .K4_C2_W1(32'hbe06a6f3), .K4_C2_W2(32'hbc9e9679), .K4_C2_W3(32'hbe29548a), .K4_C2_W4(32'h3d9b32d6), .K4_C2_W5(32'h3cbec723), .K4_C2_W6(32'h3dc8a60b), .K4_C2_W7(32'h3d3f55b2), .K4_C2_W8(32'hbd0876b3), 
		.K4_C3_W0(32'hbcb6e5b8), .K4_C3_W1(32'h3d4e1d11), .K4_C3_W2(32'hbd8906be), .K4_C3_W3(32'hbe29a530), .K4_C3_W4(32'hbde3c274), .K4_C3_W5(32'hbd562a58), .K4_C3_W6(32'hbd15ee4a), .K4_C3_W7(32'h3ce60be9), .K4_C3_W8(32'h3d1021e3), 
		.K4_C4_W0(32'hbdacce25), .K4_C4_W1(32'hbdeb2080), .K4_C4_W2(32'h3bdfc4a2), .K4_C4_W3(32'h3e2bd93d), .K4_C4_W4(32'h3ca5252f), .K4_C4_W5(32'hbdc7526c), .K4_C4_W6(32'hbd6c605f), .K4_C4_W7(32'h3daae1a2), .K4_C4_W8(32'hbbfbb6e4), 
		.K4_C5_W0(32'h3d82a20a), .K4_C5_W1(32'h3e0579e4), .K4_C5_W2(32'hbdc59e00), .K4_C5_W3(32'hbe13bbbe), .K4_C5_W4(32'hbc475c1d), .K4_C5_W5(32'h3dd6b23f), .K4_C5_W6(32'hbb2f5cd2), .K4_C5_W7(32'h3d4daa95), .K4_C5_W8(32'h3cd3460c), 
		.K4_C6_W0(32'h3ded104f), .K4_C6_W1(32'h3b90771a), .K4_C6_W2(32'hbdc9dde8), .K4_C6_W3(32'hbdb2f167), .K4_C6_W4(32'h3d445e8d), .K4_C6_W5(32'hbdee3994), .K4_C6_W6(32'hbc7d80af), .K4_C6_W7(32'hbdaff768), .K4_C6_W8(32'h3d21570e), 
		.K4_C7_W0(32'h3df17767), .K4_C7_W1(32'hbd07add9), .K4_C7_W2(32'hbe16ca40), .K4_C7_W3(32'h3d581921), .K4_C7_W4(32'hbe218891), .K4_C7_W5(32'hbe0451d0), .K4_C7_W6(32'h3e0011af), .K4_C7_W7(32'h3d99ce4d), .K4_C7_W8(32'hbd076f15), 
		.K4_C8_W0(32'h3d5ff3bc), .K4_C8_W1(32'hba86f81b), .K4_C8_W2(32'h3ca6a695), .K4_C8_W3(32'h3d9c320a), .K4_C8_W4(32'h3df03b25), .K4_C8_W5(32'h3e02086e), .K4_C8_W6(32'h3c992e72), .K4_C8_W7(32'h3d9091d5), .K4_C8_W8(32'h3da2ced6), 
		.K4_C9_W0(32'h3c8d001f), .K4_C9_W1(32'h3e25fae1), .K4_C9_W2(32'hbcd78bda), .K4_C9_W3(32'h3d6c5723), .K4_C9_W4(32'h3dc01c98), .K4_C9_W5(32'hbd9c4923), .K4_C9_W6(32'h3dc7fda5), .K4_C9_W7(32'hbd9bf777), .K4_C9_W8(32'hbe0079b3), 
		.K4_C10_W0(32'h3d88d552), .K4_C10_W1(32'h3d5a05ba), .K4_C10_W2(32'hbd4f368f), .K4_C10_W3(32'hbe14bc55), .K4_C10_W4(32'hbe1abe01), .K4_C10_W5(32'h3dae144f), .K4_C10_W6(32'h3e2a7cf5), .K4_C10_W7(32'hbc7f80bb), .K4_C10_W8(32'h3e01a981), 
		.K4_C11_W0(32'h3cc9ccb3), .K4_C11_W1(32'hbd9391af), .K4_C11_W2(32'h3ac00471), .K4_C11_W3(32'hbe0ec218), .K4_C11_W4(32'h3dbc75a7), .K4_C11_W5(32'hbe014438), .K4_C11_W6(32'hbd715387), .K4_C11_W7(32'h3e15436f), .K4_C11_W8(32'h3e129f4f), 
		.K4_C12_W0(32'hbdcb17c0), .K4_C12_W1(32'h3d3fa84f), .K4_C12_W2(32'hbd5392c5), .K4_C12_W3(32'hbd32bbfc), .K4_C12_W4(32'hbd502271), .K4_C12_W5(32'h3db6b1c3), .K4_C12_W6(32'hbd93f893), .K4_C12_W7(32'h3d664c55), .K4_C12_W8(32'hbcbc34da), 
		.K4_C13_W0(32'hbd63ac45), .K4_C13_W1(32'hbdfe9351), .K4_C13_W2(32'h3cb4985e), .K4_C13_W3(32'h3dd3b801), .K4_C13_W4(32'hbddd65dc), .K4_C13_W5(32'hbdde5d0a), .K4_C13_W6(32'hbd6e701e), .K4_C13_W7(32'h3cf628dd), .K4_C13_W8(32'hbde333e3), 
		.K4_C14_W0(32'h3d88a794), .K4_C14_W1(32'h3d5cc404), .K4_C14_W2(32'hbd376a3a), .K4_C14_W3(32'hbdf656c1), .K4_C14_W4(32'hbd3ca266), .K4_C14_W5(32'hbc972b86), .K4_C14_W6(32'hbdd95e6c), .K4_C14_W7(32'hbd32edf9), .K4_C14_W8(32'hbdb12e3c), 
		.K4_C15_W0(32'hbd07cbd3), .K4_C15_W1(32'h3dfb7542), .K4_C15_W2(32'h3dba6f65), .K4_C15_W3(32'h3cca82e5), .K4_C15_W4(32'h3dc77f97), .K4_C15_W5(32'h3e07cc66), .K4_C15_W6(32'hbd8db882), .K4_C15_W7(32'hbd1f8f85), .K4_C15_W8(32'h3dc7a365), 
		.K4_BIAS (32'h3d0bb565),

		.K5_C0_W0(32'hbcd4d670), .K5_C0_W1(32'hbca733f9), .K5_C0_W2(32'h3dd21987), .K5_C0_W3(32'h3ca295dc), .K5_C0_W4(32'h3e2152ad), .K5_C0_W5(32'h3d990668), .K5_C0_W6(32'h3c5c7783), .K5_C0_W7(32'h3d923fc5), .K5_C0_W8(32'hbb8ab223), 
		.K5_C1_W0(32'h3d038300), .K5_C1_W1(32'hbe013724), .K5_C1_W2(32'hbdf2619a), .K5_C1_W3(32'hbda92110), .K5_C1_W4(32'hbd19078c), .K5_C1_W5(32'hbdbf0ef1), .K5_C1_W6(32'hbe0cdb9a), .K5_C1_W7(32'hbd63fb29), .K5_C1_W8(32'h3d3ce419), 
		.K5_C2_W0(32'hbdb25f9c), .K5_C2_W1(32'h3dc55cd6), .K5_C2_W2(32'hbd1f4d6b), .K5_C2_W3(32'hbe07af62), .K5_C2_W4(32'h3d536414), .K5_C2_W5(32'hbd8bbd79), .K5_C2_W6(32'h3e05a12d), .K5_C2_W7(32'hbe02313f), .K5_C2_W8(32'h3cf147cf), 
		.K5_C3_W0(32'hbcdb9be4), .K5_C3_W1(32'h3dd7796c), .K5_C3_W2(32'hbe185f43), .K5_C3_W3(32'hbdb11456), .K5_C3_W4(32'h3dba7da9), .K5_C3_W5(32'h3d2b7873), .K5_C3_W6(32'hbd4562b1), .K5_C3_W7(32'h3d4ecbaf), .K5_C3_W8(32'hbe113863), 
		.K5_C4_W0(32'h3d40f2f4), .K5_C4_W1(32'hbd4bb08f), .K5_C4_W2(32'hbd842a9f), .K5_C4_W3(32'hbc09a606), .K5_C4_W4(32'h3cdcc5a8), .K5_C4_W5(32'h3d0300f7), .K5_C4_W6(32'h3d59ed98), .K5_C4_W7(32'hbba69239), .K5_C4_W8(32'h3e096602), 
		.K5_C5_W0(32'hbe1b48a1), .K5_C5_W1(32'hbb65b7f0), .K5_C5_W2(32'h3da06c09), .K5_C5_W3(32'hbe22165a), .K5_C5_W4(32'hbb1470f0), .K5_C5_W5(32'h3d375d8d), .K5_C5_W6(32'h3e14a1fe), .K5_C5_W7(32'h3be04926), .K5_C5_W8(32'hbb3590a5), 
		.K5_C6_W0(32'h3cc9324c), .K5_C6_W1(32'hbdae145c), .K5_C6_W2(32'hbd6905f8), .K5_C6_W3(32'h3d91f2f4), .K5_C6_W4(32'hbd5f0e8b), .K5_C6_W5(32'h3d5b483f), .K5_C6_W6(32'hbd2b5074), .K5_C6_W7(32'h3a30c7ca), .K5_C6_W8(32'hbb97778c), 
		.K5_C7_W0(32'hbcf35c6c), .K5_C7_W1(32'hbc51680f), .K5_C7_W2(32'h3d4ca4e6), .K5_C7_W3(32'h3dd4a7a9), .K5_C7_W4(32'hbddeb16a), .K5_C7_W5(32'hbab2086a), .K5_C7_W6(32'h3dcee96a), .K5_C7_W7(32'h3da14e05), .K5_C7_W8(32'hbd4f120e), 
		.K5_C8_W0(32'h3dbab65b), .K5_C8_W1(32'hbce53330), .K5_C8_W2(32'h3db0e823), .K5_C8_W3(32'h3d4eb43d), .K5_C8_W4(32'h3c0b0e3f), .K5_C8_W5(32'h3d386bf5), .K5_C8_W6(32'h3d9ff4f4), .K5_C8_W7(32'hbcfc547c), .K5_C8_W8(32'hbd0c388a), 
		.K5_C9_W0(32'hbdb8315b), .K5_C9_W1(32'hbd91ddac), .K5_C9_W2(32'hbdd2d7c2), .K5_C9_W3(32'h3d214e7a), .K5_C9_W4(32'hbdb89409), .K5_C9_W5(32'hbe1f2793), .K5_C9_W6(32'hbd57c6c1), .K5_C9_W7(32'hbc0cb252), .K5_C9_W8(32'h3e206a3f), 
		.K5_C10_W0(32'hbdb4de0a), .K5_C10_W1(32'hbda2fcad), .K5_C10_W2(32'h3e20a44d), .K5_C10_W3(32'hbda5bd1e), .K5_C10_W4(32'h3e0753fe), .K5_C10_W5(32'h3e08970a), .K5_C10_W6(32'hbc8bc505), .K5_C10_W7(32'hbbf4b3c6), .K5_C10_W8(32'hbd854a1a), 
		.K5_C11_W0(32'hbdcf614a), .K5_C11_W1(32'hbd2e4002), .K5_C11_W2(32'hbc248fbf), .K5_C11_W3(32'h3e05245a), .K5_C11_W4(32'h3e125c8e), .K5_C11_W5(32'hbdd5dd1e), .K5_C11_W6(32'h3dfbd86c), .K5_C11_W7(32'hbb908acc), .K5_C11_W8(32'hbde18159), 
		.K5_C12_W0(32'h3e2d4bf8), .K5_C12_W1(32'h3e0a1238), .K5_C12_W2(32'hbbbb750a), .K5_C12_W3(32'h3dee5982), .K5_C12_W4(32'h3d7d426c), .K5_C12_W5(32'hbe057aaf), .K5_C12_W6(32'h3b3f4cfb), .K5_C12_W7(32'h3d917512), .K5_C12_W8(32'hbda2c448), 
		.K5_C13_W0(32'h3d190e04), .K5_C13_W1(32'hbc7cd4cd), .K5_C13_W2(32'hbde14032), .K5_C13_W3(32'hbcdb9ae8), .K5_C13_W4(32'hbe40adc8), .K5_C13_W5(32'h3cf7b2e5), .K5_C13_W6(32'hbd1de366), .K5_C13_W7(32'h3da5baeb), .K5_C13_W8(32'h3e122d8d), 
		.K5_C14_W0(32'h3c83b7d2), .K5_C14_W1(32'h3ce5a47b), .K5_C14_W2(32'h3d9ba9f4), .K5_C14_W3(32'hbded9a1d), .K5_C14_W4(32'h3e05bec3), .K5_C14_W5(32'h3d0e08b5), .K5_C14_W6(32'h3d1bface), .K5_C14_W7(32'h3c62a677), .K5_C14_W8(32'hbe075c08), 
		.K5_C15_W0(32'h3d644d47), .K5_C15_W1(32'h3ca817ec), .K5_C15_W2(32'h3b2caec6), .K5_C15_W3(32'hbe0d9f82), .K5_C15_W4(32'h3d7fe009), .K5_C15_W5(32'hbd8afdec), .K5_C15_W6(32'hbe251771), .K5_C15_W7(32'h3d60983e), .K5_C15_W8(32'hbd106445), 
		.K5_BIAS (32'h3ce4caf4),

		.K6_C0_W0(32'h3d19d22e), .K6_C0_W1(32'hbc62af15), .K6_C0_W2(32'h3d65f44e), .K6_C0_W3(32'h3d08a573), .K6_C0_W4(32'h3bab2254), .K6_C0_W5(32'h3dbaa57d), .K6_C0_W6(32'h3de42379), .K6_C0_W7(32'h3da5117b), .K6_C0_W8(32'h3e02f78a), 
		.K6_C1_W0(32'hbdf8c588), .K6_C1_W1(32'h3db9c1f7), .K6_C1_W2(32'h3c852583), .K6_C1_W3(32'h3db35cfc), .K6_C1_W4(32'hbd5ddbbb), .K6_C1_W5(32'hbde5f5ee), .K6_C1_W6(32'h3daf172e), .K6_C1_W7(32'hbe017375), .K6_C1_W8(32'h3d053d5c), 
		.K6_C2_W0(32'h3dbc23cc), .K6_C2_W1(32'hbdbc71f0), .K6_C2_W2(32'h3cac81c0), .K6_C2_W3(32'hbe036580), .K6_C2_W4(32'hbe2a203b), .K6_C2_W5(32'hbdb0ef7e), .K6_C2_W6(32'h3ddce25e), .K6_C2_W7(32'h3da1bd22), .K6_C2_W8(32'h3d66fa93), 
		.K6_C3_W0(32'h3d5d801b), .K6_C3_W1(32'h3dde0e84), .K6_C3_W2(32'hbddd5f5f), .K6_C3_W3(32'hbe0684c8), .K6_C3_W4(32'h3dfac2a4), .K6_C3_W5(32'h3a5c5d14), .K6_C3_W6(32'hbdafdc17), .K6_C3_W7(32'hbe12d9f2), .K6_C3_W8(32'hbd37b007), 
		.K6_C4_W0(32'h3e2d4669), .K6_C4_W1(32'hbd1088a9), .K6_C4_W2(32'h3e281d4c), .K6_C4_W3(32'h3d53aff7), .K6_C4_W4(32'h3e2bc373), .K6_C4_W5(32'h3dd09754), .K6_C4_W6(32'hbdb101cb), .K6_C4_W7(32'h3df05cc5), .K6_C4_W8(32'h3d707b14), 
		.K6_C5_W0(32'hbd013ca7), .K6_C5_W1(32'h3c111d8d), .K6_C5_W2(32'hbda296ee), .K6_C5_W3(32'hbd183a1c), .K6_C5_W4(32'hbe0e744c), .K6_C5_W5(32'hbde7108a), .K6_C5_W6(32'hbdd9551d), .K6_C5_W7(32'h3d61838d), .K6_C5_W8(32'h3e0adeaf), 
		.K6_C6_W0(32'h3e11b449), .K6_C6_W1(32'h3d8a4fd3), .K6_C6_W2(32'hbd102ea1), .K6_C6_W3(32'h3c9df94b), .K6_C6_W4(32'hba84dcc6), .K6_C6_W5(32'h3d6ae203), .K6_C6_W6(32'h3d1c01eb), .K6_C6_W7(32'h3db9973f), .K6_C6_W8(32'hbdc86636), 
		.K6_C7_W0(32'h3d00ee1e), .K6_C7_W1(32'hbd80ea73), .K6_C7_W2(32'hbdcd1f97), .K6_C7_W3(32'hbd39b797), .K6_C7_W4(32'hbd3518f3), .K6_C7_W5(32'h3d158d2a), .K6_C7_W6(32'hbda2ac9b), .K6_C7_W7(32'hbd0ebed5), .K6_C7_W8(32'hbd8c2e17), 
		.K6_C8_W0(32'hbe533ff5), .K6_C8_W1(32'hbe48dc6c), .K6_C8_W2(32'hbe018252), .K6_C8_W3(32'h3b56bdc3), .K6_C8_W4(32'hbcbd286a), .K6_C8_W5(32'hbd9dba1a), .K6_C8_W6(32'h3df35d3e), .K6_C8_W7(32'hbdc45b65), .K6_C8_W8(32'hbd955604), 
		.K6_C9_W0(32'h3d9f9662), .K6_C9_W1(32'h3bfd830f), .K6_C9_W2(32'h3db00597), .K6_C9_W3(32'h3df6f986), .K6_C9_W4(32'h3e21ffec), .K6_C9_W5(32'h3e1acf64), .K6_C9_W6(32'hbd88169c), .K6_C9_W7(32'h3dd2752e), .K6_C9_W8(32'h3d9802b2), 
		.K6_C10_W0(32'h3de37d1a), .K6_C10_W1(32'h3dcc768f), .K6_C10_W2(32'hbe2d6a5f), .K6_C10_W3(32'hbdcfa32d), .K6_C10_W4(32'h3da8b119), .K6_C10_W5(32'hbc66a141), .K6_C10_W6(32'hbd599842), .K6_C10_W7(32'h3db9d191), .K6_C10_W8(32'h3da3f220), 
		.K6_C11_W0(32'hbd445087), .K6_C11_W1(32'h3c9d6dc5), .K6_C11_W2(32'h3d1e64cc), .K6_C11_W3(32'h3d266ed1), .K6_C11_W4(32'h3df54ec0), .K6_C11_W5(32'hbdba840f), .K6_C11_W6(32'hbde64b82), .K6_C11_W7(32'hbd3ffca0), .K6_C11_W8(32'h3db6b1bd), 
		.K6_C12_W0(32'h3cfa879a), .K6_C12_W1(32'h3d4f385b), .K6_C12_W2(32'hbd380510), .K6_C12_W3(32'hbd107153), .K6_C12_W4(32'h3dea6dca), .K6_C12_W5(32'hbe1339cf), .K6_C12_W6(32'h3d3d760a), .K6_C12_W7(32'h3dfad915), .K6_C12_W8(32'h3d52bc3d), 
		.K6_C13_W0(32'h3e314121), .K6_C13_W1(32'h3dc8b6cb), .K6_C13_W2(32'h3d3de626), .K6_C13_W3(32'h3d5d35b8), .K6_C13_W4(32'h3e155cba), .K6_C13_W5(32'h3d23e9b8), .K6_C13_W6(32'h3d82cf3c), .K6_C13_W7(32'hbe026130), .K6_C13_W8(32'hbd054400), 
		.K6_C14_W0(32'hbe1d51c1), .K6_C14_W1(32'h3cf188d1), .K6_C14_W2(32'hbcaf9909), .K6_C14_W3(32'h3d8da024), .K6_C14_W4(32'h3b788349), .K6_C14_W5(32'h3d928202), .K6_C14_W6(32'hbe00e46c), .K6_C14_W7(32'h3daca73e), .K6_C14_W8(32'h3d566e44), 
		.K6_C15_W0(32'h3c894c72), .K6_C15_W1(32'hbd9c01ac), .K6_C15_W2(32'hbdc03683), .K6_C15_W3(32'hbd732141), .K6_C15_W4(32'h3d410419), .K6_C15_W5(32'hbd82af68), .K6_C15_W6(32'hbd84301a), .K6_C15_W7(32'h3d5a172f), .K6_C15_W8(32'h3d736243), 
		.K6_BIAS (32'h3d86eb4b),

		.K7_C0_W0(32'h3cacbf35), .K7_C0_W1(32'hbe07d5c7), .K7_C0_W2(32'h3d659ec9), .K7_C0_W3(32'hbc8a181b), .K7_C0_W4(32'hbe0b7a11), .K7_C0_W5(32'hbdc814bc), .K7_C0_W6(32'hbe07cc9b), .K7_C0_W7(32'h3d55f059), .K7_C0_W8(32'h3bc5b2a2), 
		.K7_C1_W0(32'h3da241cc), .K7_C1_W1(32'hbd948f3c), .K7_C1_W2(32'h3e0913da), .K7_C1_W3(32'h3cb19644), .K7_C1_W4(32'h3da7d76a), .K7_C1_W5(32'h3b3cf176), .K7_C1_W6(32'h3bd60367), .K7_C1_W7(32'h3df2bdef), .K7_C1_W8(32'hbe193169), 
		.K7_C2_W0(32'hbdcb30b3), .K7_C2_W1(32'h3db90b36), .K7_C2_W2(32'hbe07de65), .K7_C2_W3(32'h3d4794a8), .K7_C2_W4(32'h3d1dbf3b), .K7_C2_W5(32'h3e0601c1), .K7_C2_W6(32'hbd7a93bc), .K7_C2_W7(32'hbdbeeecf), .K7_C2_W8(32'hbdfd2bdb), 
		.K7_C3_W0(32'hbe32de8a), .K7_C3_W1(32'h3e142b79), .K7_C3_W2(32'h3e07810a), .K7_C3_W3(32'hbe1b6e85), .K7_C3_W4(32'h3aa835a9), .K7_C3_W5(32'hbe28e55f), .K7_C3_W6(32'hbd50fc4d), .K7_C3_W7(32'hbced2066), .K7_C3_W8(32'h3e3414a6), 
		.K7_C4_W0(32'h3c22a998), .K7_C4_W1(32'hbccc100c), .K7_C4_W2(32'h3d6c7f6e), .K7_C4_W3(32'h3e00781a), .K7_C4_W4(32'h3e337c61), .K7_C4_W5(32'h3dd357cb), .K7_C4_W6(32'h39fb52ba), .K7_C4_W7(32'h3dc0311e), .K7_C4_W8(32'h3dd2ecaf), 
		.K7_C5_W0(32'h3b759ce5), .K7_C5_W1(32'hbcf3dbab), .K7_C5_W2(32'h3dd8b230), .K7_C5_W3(32'h3d95fd76), .K7_C5_W4(32'h3e4085a3), .K7_C5_W5(32'h3c6ff11e), .K7_C5_W6(32'hbbfc8a1e), .K7_C5_W7(32'h3dd9ad58), .K7_C5_W8(32'hbd290fa7), 
		.K7_C6_W0(32'hbdd97c39), .K7_C6_W1(32'h3c97306c), .K7_C6_W2(32'h3d47afb4), .K7_C6_W3(32'h3ce41dd6), .K7_C6_W4(32'hbd47ba07), .K7_C6_W5(32'h3d181e64), .K7_C6_W6(32'hbe01ed63), .K7_C6_W7(32'h3da5b519), .K7_C6_W8(32'h3c2be34a), 
		.K7_C7_W0(32'h3debd273), .K7_C7_W1(32'h3a941682), .K7_C7_W2(32'h3d49229d), .K7_C7_W3(32'hbc91ca82), .K7_C7_W4(32'hbba43e9d), .K7_C7_W5(32'h3dc94bfb), .K7_C7_W6(32'h3d218555), .K7_C7_W7(32'h3dc6d793), .K7_C7_W8(32'h3d759341), 
		.K7_C8_W0(32'h3de46450), .K7_C8_W1(32'hbe20bc90), .K7_C8_W2(32'hbc8d8776), .K7_C8_W3(32'hbe0c3224), .K7_C8_W4(32'hbdb43e89), .K7_C8_W5(32'h3d1e53ce), .K7_C8_W6(32'hbd822f6c), .K7_C8_W7(32'hbdac248e), .K7_C8_W8(32'h3b498904), 
		.K7_C9_W0(32'h3e14f43b), .K7_C9_W1(32'h3d877c42), .K7_C9_W2(32'hbd429e8e), .K7_C9_W3(32'h3e28a4b8), .K7_C9_W4(32'h3e3840f7), .K7_C9_W5(32'h3dbc10ea), .K7_C9_W6(32'hbc93080f), .K7_C9_W7(32'hba7a4075), .K7_C9_W8(32'hbe08a9bc), 
		.K7_C10_W0(32'hbd08b886), .K7_C10_W1(32'h3e1a9356), .K7_C10_W2(32'hbdc60909), .K7_C10_W3(32'h3dd552f1), .K7_C10_W4(32'h3d935f0c), .K7_C10_W5(32'h3dcc3f7d), .K7_C10_W6(32'h3d8b1631), .K7_C10_W7(32'hbe011461), .K7_C10_W8(32'hbd6a81bb), 
		.K7_C11_W0(32'hbd1a538e), .K7_C11_W1(32'hbe06ed1b), .K7_C11_W2(32'hbdd5da8d), .K7_C11_W3(32'hbde6038e), .K7_C11_W4(32'hbe22b9b8), .K7_C11_W5(32'hbe0d14d6), .K7_C11_W6(32'h3e0ba0db), .K7_C11_W7(32'hbd9185eb), .K7_C11_W8(32'h3deaf539), 
		.K7_C12_W0(32'hbbc7de53), .K7_C12_W1(32'hbd6f0c46), .K7_C12_W2(32'h3c030665), .K7_C12_W3(32'h3d0a4376), .K7_C12_W4(32'hbdb65e44), .K7_C12_W5(32'h3cfb7aef), .K7_C12_W6(32'h3dc8cbb7), .K7_C12_W7(32'h3bef0922), .K7_C12_W8(32'h3cb456ab), 
		.K7_C13_W0(32'h3e0c327a), .K7_C13_W1(32'h3def3292), .K7_C13_W2(32'h3dcec7eb), .K7_C13_W3(32'h3ca7d221), .K7_C13_W4(32'h3e2b01fd), .K7_C13_W5(32'hbc119888), .K7_C13_W6(32'hbd7670f6), .K7_C13_W7(32'hbd926017), .K7_C13_W8(32'hbdf5f4fe), 
		.K7_C14_W0(32'h3dae1054), .K7_C14_W1(32'hbd860d3c), .K7_C14_W2(32'hbcc428e1), .K7_C14_W3(32'hbdf30632), .K7_C14_W4(32'h3ccb1d50), .K7_C14_W5(32'hbb44025f), .K7_C14_W6(32'h3b99c4dc), .K7_C14_W7(32'h3d854d82), .K7_C14_W8(32'h3e2d78c2), 
		.K7_C15_W0(32'h3dd7f3ce), .K7_C15_W1(32'h3dc121a4), .K7_C15_W2(32'hbd61433b), .K7_C15_W3(32'h3d2c649f), .K7_C15_W4(32'h3b1b8dbb), .K7_C15_W5(32'h3dfb505c), .K7_C15_W6(32'hbe054e69), .K7_C15_W7(32'h3e041ef7), .K7_C15_W8(32'h3e1088b7), 
		.K7_BIAS (32'hbb17a59c),

		.K8_C0_W0(32'hbd064f3d), .K8_C0_W1(32'h3cdb21cd), .K8_C0_W2(32'h3d2a1bb4), .K8_C0_W3(32'h3d44990b), .K8_C0_W4(32'hbcd2f40e), .K8_C0_W5(32'h3d926772), .K8_C0_W6(32'h3d823c16), .K8_C0_W7(32'h3da020d8), .K8_C0_W8(32'h3a5e7b8e), 
		.K8_C1_W0(32'h3b1b802d), .K8_C1_W1(32'h3d6dd130), .K8_C1_W2(32'hbce62fad), .K8_C1_W3(32'h3dc8ddb1), .K8_C1_W4(32'hbdd74e0f), .K8_C1_W5(32'h3d8b38e5), .K8_C1_W6(32'h3d0c25c7), .K8_C1_W7(32'hbdd82af3), .K8_C1_W8(32'hbd4fbe2b), 
		.K8_C2_W0(32'hbdce4922), .K8_C2_W1(32'h3e1ce2aa), .K8_C2_W2(32'h3d3016b4), .K8_C2_W3(32'h3c428071), .K8_C2_W4(32'h3d09991e), .K8_C2_W5(32'h3dd6548f), .K8_C2_W6(32'hbdb92d4c), .K8_C2_W7(32'hbd914340), .K8_C2_W8(32'hbdce3a5d), 
		.K8_C3_W0(32'h3d26e010), .K8_C3_W1(32'hbdc2c3ff), .K8_C3_W2(32'h3d8b7dff), .K8_C3_W3(32'hbda16fc4), .K8_C3_W4(32'h3df19a3b), .K8_C3_W5(32'h3e099053), .K8_C3_W6(32'hbde4ee51), .K8_C3_W7(32'h3d84ea8f), .K8_C3_W8(32'h3e22e889), 
		.K8_C4_W0(32'h3c52f8cf), .K8_C4_W1(32'h3ceeca44), .K8_C4_W2(32'h3d807a0b), .K8_C4_W3(32'hbdaa84a6), .K8_C4_W4(32'hbc72ea55), .K8_C4_W5(32'h3dca5835), .K8_C4_W6(32'h3d4b297e), .K8_C4_W7(32'hbe021285), .K8_C4_W8(32'hbdfd3c72), 
		.K8_C5_W0(32'hbc329b74), .K8_C5_W1(32'h3e081c3f), .K8_C5_W2(32'h3e18d47c), .K8_C5_W3(32'hbe010c40), .K8_C5_W4(32'hbe1c5421), .K8_C5_W5(32'hbb5b255c), .K8_C5_W6(32'h3d9db93f), .K8_C5_W7(32'h3ba09ea9), .K8_C5_W8(32'hbd4511b5), 
		.K8_C6_W0(32'h3e0ecfc2), .K8_C6_W1(32'hbda95b54), .K8_C6_W2(32'h3e26daf3), .K8_C6_W3(32'hbd2cc68c), .K8_C6_W4(32'hbd3d9c70), .K8_C6_W5(32'hbd8840b7), .K8_C6_W6(32'h3e11e728), .K8_C6_W7(32'hbdf523b9), .K8_C6_W8(32'h3af9529a), 
		.K8_C7_W0(32'hbd81e19c), .K8_C7_W1(32'hbdf91e61), .K8_C7_W2(32'h3d6963ec), .K8_C7_W3(32'hbc413906), .K8_C7_W4(32'hbd2e0f9d), .K8_C7_W5(32'hbe078662), .K8_C7_W6(32'hbdf6ac6a), .K8_C7_W7(32'hbe1d0e31), .K8_C7_W8(32'hbd85e578), 
		.K8_C8_W0(32'hbca5c4db), .K8_C8_W1(32'h3d0559f4), .K8_C8_W2(32'h3d232983), .K8_C8_W3(32'hbcee5970), .K8_C8_W4(32'hbd8b7a0c), .K8_C8_W5(32'hbdbc80e2), .K8_C8_W6(32'h3de45e99), .K8_C8_W7(32'hbd13093b), .K8_C8_W8(32'h3dd180c9), 
		.K8_C9_W0(32'h3d79c0e2), .K8_C9_W1(32'h3e0e573f), .K8_C9_W2(32'hbcdab1f6), .K8_C9_W3(32'hbe073146), .K8_C9_W4(32'h3dcbd2d5), .K8_C9_W5(32'hbe005102), .K8_C9_W6(32'hbd0f1cad), .K8_C9_W7(32'hbdfa3618), .K8_C9_W8(32'h3d820ab1), 
		.K8_C10_W0(32'h3df2022e), .K8_C10_W1(32'h3d762aaa), .K8_C10_W2(32'h3d9b62e5), .K8_C10_W3(32'hbde9d0d1), .K8_C10_W4(32'hba1a1285), .K8_C10_W5(32'hbda32438), .K8_C10_W6(32'h3da522f0), .K8_C10_W7(32'h3db7bba0), .K8_C10_W8(32'hbe25774c), 
		.K8_C11_W0(32'hbd969ce0), .K8_C11_W1(32'h3b967cf3), .K8_C11_W2(32'hbbdc9226), .K8_C11_W3(32'h3d2e02ac), .K8_C11_W4(32'h3e1c8315), .K8_C11_W5(32'hbab1f9fa), .K8_C11_W6(32'h3c87f834), .K8_C11_W7(32'hbdcacdef), .K8_C11_W8(32'h3dc7999a), 
		.K8_C12_W0(32'h3d6cdbd9), .K8_C12_W1(32'h3de8533e), .K8_C12_W2(32'h3d3c5ed2), .K8_C12_W3(32'h3da9e90d), .K8_C12_W4(32'hbe05aa0a), .K8_C12_W5(32'hbc67c692), .K8_C12_W6(32'hbcfae6e5), .K8_C12_W7(32'h3de38e7d), .K8_C12_W8(32'h3c66f2cd), 
		.K8_C13_W0(32'h3d94954e), .K8_C13_W1(32'h3d156685), .K8_C13_W2(32'h3d8633cb), .K8_C13_W3(32'h3e0057b8), .K8_C13_W4(32'hbdf99321), .K8_C13_W5(32'hbdc9ec1e), .K8_C13_W6(32'hbc8f4564), .K8_C13_W7(32'hbdf05d92), .K8_C13_W8(32'hbdc8a7f9), 
		.K8_C14_W0(32'hbdc63211), .K8_C14_W1(32'hbdf207ac), .K8_C14_W2(32'h3cd8ac21), .K8_C14_W3(32'hbdf3bace), .K8_C14_W4(32'h3e07cafc), .K8_C14_W5(32'hbe036d78), .K8_C14_W6(32'hbd2835be), .K8_C14_W7(32'h3e06131e), .K8_C14_W8(32'h3ded1a99), 
		.K8_C15_W0(32'h3c9d4d65), .K8_C15_W1(32'h3dfbe7c2), .K8_C15_W2(32'hbda82190), .K8_C15_W3(32'h3da23205), .K8_C15_W4(32'h3d943a03), .K8_C15_W5(32'hbd6fbcda), .K8_C15_W6(32'h3cf87df2), .K8_C15_W7(32'hbd501cb5), .K8_C15_W8(32'h3da6407a), 
		.K8_BIAS (32'hbcb94f4f),

		.K9_C0_W0(32'hbcd907c8), .K9_C0_W1(32'hbdf8a2aa), .K9_C0_W2(32'hbcddb282), .K9_C0_W3(32'hbce3c558), .K9_C0_W4(32'h3d8d1aad), .K9_C0_W5(32'hbdbae14c), .K9_C0_W6(32'h3db9354f), .K9_C0_W7(32'h3e2529c0), .K9_C0_W8(32'h3d709a40), 
		.K9_C1_W0(32'hbd686f45), .K9_C1_W1(32'hbd1b40a0), .K9_C1_W2(32'hbe08e643), .K9_C1_W3(32'h3d873fa3), .K9_C1_W4(32'h3df0c1eb), .K9_C1_W5(32'h3dda436b), .K9_C1_W6(32'hbe1ddb6f), .K9_C1_W7(32'hbb3333e4), .K9_C1_W8(32'h3dc09763), 
		.K9_C2_W0(32'hbd5c9688), .K9_C2_W1(32'h3dc69073), .K9_C2_W2(32'h3e0c6857), .K9_C2_W3(32'h3dbf73e3), .K9_C2_W4(32'h3e113c20), .K9_C2_W5(32'h3c0eb12b), .K9_C2_W6(32'h3dc4c594), .K9_C2_W7(32'hbde62f22), .K9_C2_W8(32'hbbdc48dd), 
		.K9_C3_W0(32'hbc7747f5), .K9_C3_W1(32'h3dd218f4), .K9_C3_W2(32'hbdc1a5f3), .K9_C3_W3(32'h3dacd3c0), .K9_C3_W4(32'hbdab2607), .K9_C3_W5(32'hbdcc8f6b), .K9_C3_W6(32'h3e00af4d), .K9_C3_W7(32'h3d92209b), .K9_C3_W8(32'h3e06ab6d), 
		.K9_C4_W0(32'hbdca7be6), .K9_C4_W1(32'hbe188933), .K9_C4_W2(32'h3e0466e9), .K9_C4_W3(32'hbdfe4bab), .K9_C4_W4(32'hbd6b45cd), .K9_C4_W5(32'h3dacc141), .K9_C4_W6(32'hbdb5ad67), .K9_C4_W7(32'hbdb0b471), .K9_C4_W8(32'hbd4068d0), 
		.K9_C5_W0(32'h3d9db7ac), .K9_C5_W1(32'hb9ec5cc6), .K9_C5_W2(32'h3da6f445), .K9_C5_W3(32'hbc85c48d), .K9_C5_W4(32'hbdefb135), .K9_C5_W5(32'hbdddeaf5), .K9_C5_W6(32'h3df34efb), .K9_C5_W7(32'h3de0bf79), .K9_C5_W8(32'hba43aeb4), 
		.K9_C6_W0(32'h3d0c1557), .K9_C6_W1(32'h3df8b480), .K9_C6_W2(32'hbdbd38b2), .K9_C6_W3(32'h3cb4a73c), .K9_C6_W4(32'hbe2d65c6), .K9_C6_W5(32'hbd5b04b4), .K9_C6_W6(32'hbe209a0d), .K9_C6_W7(32'hbdc20d87), .K9_C6_W8(32'hbe2a8bd0), 
		.K9_C7_W0(32'hbb332dbc), .K9_C7_W1(32'hbd8116ad), .K9_C7_W2(32'h3da03711), .K9_C7_W3(32'hbd8f86f7), .K9_C7_W4(32'h3d58a2a5), .K9_C7_W5(32'hbd423edf), .K9_C7_W6(32'h3d903a12), .K9_C7_W7(32'h3d9bc81d), .K9_C7_W8(32'h3d53b7bf), 
		.K9_C8_W0(32'h3dc9be9a), .K9_C8_W1(32'h3d61fd2f), .K9_C8_W2(32'h3dc1f516), .K9_C8_W3(32'hbd56e218), .K9_C8_W4(32'h3d78787e), .K9_C8_W5(32'hbdba00d8), .K9_C8_W6(32'hbdb55f75), .K9_C8_W7(32'h3c8b269a), .K9_C8_W8(32'hbbf47016), 
		.K9_C9_W0(32'hbe12b34c), .K9_C9_W1(32'hbc420c8b), .K9_C9_W2(32'hbda02aab), .K9_C9_W3(32'hbb277fc0), .K9_C9_W4(32'hbe287cd5), .K9_C9_W5(32'h3d8d69cd), .K9_C9_W6(32'hbc3944a7), .K9_C9_W7(32'h3d812d9e), .K9_C9_W8(32'h3ddcb88a), 
		.K9_C10_W0(32'hbe086e6a), .K9_C10_W1(32'h3dec41d4), .K9_C10_W2(32'h3dfc5acd), .K9_C10_W3(32'h3dda4f55), .K9_C10_W4(32'hbd936652), .K9_C10_W5(32'hbe0736ff), .K9_C10_W6(32'hbdc84030), .K9_C10_W7(32'h3d8fbf90), .K9_C10_W8(32'hbd001371), 
		.K9_C11_W0(32'h3d08fa4f), .K9_C11_W1(32'h3da4125d), .K9_C11_W2(32'h3dde0069), .K9_C11_W3(32'hbd16be43), .K9_C11_W4(32'hbe0bf545), .K9_C11_W5(32'h3c1593f8), .K9_C11_W6(32'hbbacc368), .K9_C11_W7(32'hbceba350), .K9_C11_W8(32'hbdd129f1), 
		.K9_C12_W0(32'hbde206ae), .K9_C12_W1(32'h3dec7737), .K9_C12_W2(32'h3de10541), .K9_C12_W3(32'hbe05f22d), .K9_C12_W4(32'hbe00cb38), .K9_C12_W5(32'hbdc20873), .K9_C12_W6(32'hbd39c967), .K9_C12_W7(32'hbd72a62d), .K9_C12_W8(32'hbdd1650c), 
		.K9_C13_W0(32'hbd8a593b), .K9_C13_W1(32'h3dad11b6), .K9_C13_W2(32'h3e002e6a), .K9_C13_W3(32'hbe1541cb), .K9_C13_W4(32'h3dcc6be8), .K9_C13_W5(32'h3d74a810), .K9_C13_W6(32'hbb9cefe7), .K9_C13_W7(32'hbdcf7e92), .K9_C13_W8(32'h3d800ec4), 
		.K9_C14_W0(32'hbd74b2a6), .K9_C14_W1(32'h3df649e9), .K9_C14_W2(32'hbd8830eb), .K9_C14_W3(32'h3e0527b1), .K9_C14_W4(32'h3df07548), .K9_C14_W5(32'h3dc35c3d), .K9_C14_W6(32'h3d9ddd99), .K9_C14_W7(32'hbdd57748), .K9_C14_W8(32'hbdddee3b), 
		.K9_C15_W0(32'hbbb7983b), .K9_C15_W1(32'hbd985c90), .K9_C15_W2(32'h3df34fcc), .K9_C15_W3(32'hbcae33d9), .K9_C15_W4(32'h3c6f20d4), .K9_C15_W5(32'hbe2bf0d9), .K9_C15_W6(32'h3e0344ba), .K9_C15_W7(32'h3b139543), .K9_C15_W8(32'hbdf2c7ff), 
		.K9_BIAS (32'h3bdd4f4c),

		.K10_C0_W0(32'hbdc4231a), .K10_C0_W1(32'hbd8d2683), .K10_C0_W2(32'h3dc62da0), .K10_C0_W3(32'h3ccb1c21), .K10_C0_W4(32'hbdbac533), .K10_C0_W5(32'h3d5ea260), .K10_C0_W6(32'h3c949b03), .K10_C0_W7(32'h3e462f1d), .K10_C0_W8(32'h3cef3da3), 
		.K10_C1_W0(32'hbd0353cf), .K10_C1_W1(32'h3e157cbe), .K10_C1_W2(32'hbde49307), .K10_C1_W3(32'h3dcfae5e), .K10_C1_W4(32'h3e0f7924), .K10_C1_W5(32'hbde4c578), .K10_C1_W6(32'h3d6bfb75), .K10_C1_W7(32'h3e2d9799), .K10_C1_W8(32'h3dab75eb), 
		.K10_C2_W0(32'h3e015fd0), .K10_C2_W1(32'h3d635908), .K10_C2_W2(32'h3ca143d0), .K10_C2_W3(32'hbd576ac3), .K10_C2_W4(32'h3d0cf62d), .K10_C2_W5(32'hbe0039d3), .K10_C2_W6(32'h3d999e58), .K10_C2_W7(32'hbde5bf62), .K10_C2_W8(32'hbd99f84e), 
		.K10_C3_W0(32'hbd096378), .K10_C3_W1(32'hbdb44f37), .K10_C3_W2(32'h3c9d5cbe), .K10_C3_W3(32'h3e1f5bb0), .K10_C3_W4(32'h3d1df558), .K10_C3_W5(32'h3c80e799), .K10_C3_W6(32'hbde22fb8), .K10_C3_W7(32'hbe0cb5a4), .K10_C3_W8(32'h3d5ed38b), 
		.K10_C4_W0(32'hbde94a46), .K10_C4_W1(32'h3e10a365), .K10_C4_W2(32'hbcec303f), .K10_C4_W3(32'h3c294a7c), .K10_C4_W4(32'hbd5b833f), .K10_C4_W5(32'h3df4006a), .K10_C4_W6(32'h3e0ab67d), .K10_C4_W7(32'hbd45411b), .K10_C4_W8(32'h3d869065), 
		.K10_C5_W0(32'h3ca4bdb4), .K10_C5_W1(32'hbe0bfbe2), .K10_C5_W2(32'h3c04f30f), .K10_C5_W3(32'h3cb95efe), .K10_C5_W4(32'hbdcb27ea), .K10_C5_W5(32'hb93560c8), .K10_C5_W6(32'h3dd37f9b), .K10_C5_W7(32'hbe00767a), .K10_C5_W8(32'hbe053271), 
		.K10_C6_W0(32'hbdffa95a), .K10_C6_W1(32'h3dd61640), .K10_C6_W2(32'h3cdd91bd), .K10_C6_W3(32'hbe3a6f67), .K10_C6_W4(32'h3d1cbc71), .K10_C6_W5(32'h3dcd6c24), .K10_C6_W6(32'hbdacdc07), .K10_C6_W7(32'hbdd5cd54), .K10_C6_W8(32'h3cb2e11f), 
		.K10_C7_W0(32'h3df62165), .K10_C7_W1(32'h3d93fdfd), .K10_C7_W2(32'h3d3525d8), .K10_C7_W3(32'hbd68fb7c), .K10_C7_W4(32'h3d00924e), .K10_C7_W5(32'hbdcc718b), .K10_C7_W6(32'hbd5483fc), .K10_C7_W7(32'hbddd8deb), .K10_C7_W8(32'hbddd0430), 
		.K10_C8_W0(32'h3d145d00), .K10_C8_W1(32'h3d139485), .K10_C8_W2(32'h3de963ff), .K10_C8_W3(32'h3c0ed339), .K10_C8_W4(32'h3df57c94), .K10_C8_W5(32'h3d858af9), .K10_C8_W6(32'h3df3a57a), .K10_C8_W7(32'hbda0513f), .K10_C8_W8(32'hbcf7ff10), 
		.K10_C9_W0(32'hbd942ed3), .K10_C9_W1(32'hbdc28e43), .K10_C9_W2(32'h3dc5c75e), .K10_C9_W3(32'h3d25937d), .K10_C9_W4(32'hbd1cdf9a), .K10_C9_W5(32'h3e0ba65c), .K10_C9_W6(32'h3d50d878), .K10_C9_W7(32'hbdbb400a), .K10_C9_W8(32'h3de585a0), 
		.K10_C10_W0(32'h3d823b7d), .K10_C10_W1(32'h3df71638), .K10_C10_W2(32'hbd10f669), .K10_C10_W3(32'hbd66681f), .K10_C10_W4(32'hbdef8c48), .K10_C10_W5(32'hbdf1b6e2), .K10_C10_W6(32'hbb5c4e74), .K10_C10_W7(32'hbc8b4419), .K10_C10_W8(32'h3d8a6575), 
		.K10_C11_W0(32'h3db39b40), .K10_C11_W1(32'hbdbb7f31), .K10_C11_W2(32'hbb5b8042), .K10_C11_W3(32'hbdf1cb0e), .K10_C11_W4(32'h3948aec0), .K10_C11_W5(32'hbde31517), .K10_C11_W6(32'h3d18afdc), .K10_C11_W7(32'hbe1bae38), .K10_C11_W8(32'h3cb9f30b), 
		.K10_C12_W0(32'hbdd52e3a), .K10_C12_W1(32'h3d421e86), .K10_C12_W2(32'h3dc0ec3c), .K10_C12_W3(32'hbcf8e46d), .K10_C12_W4(32'hbccedca4), .K10_C12_W5(32'hbd76e685), .K10_C12_W6(32'h3e30cba7), .K10_C12_W7(32'h3dcc4351), .K10_C12_W8(32'h3e093ab2), 
		.K10_C13_W0(32'hbdc1fa35), .K10_C13_W1(32'h3d2e9348), .K10_C13_W2(32'h3e05303b), .K10_C13_W3(32'h3d88e61e), .K10_C13_W4(32'hbc2bec6a), .K10_C13_W5(32'h3decaaf7), .K10_C13_W6(32'h3df85337), .K10_C13_W7(32'hbcbc1ce2), .K10_C13_W8(32'h3e2873c6), 
		.K10_C14_W0(32'h3ca3eb8d), .K10_C14_W1(32'hbb1690b4), .K10_C14_W2(32'hbcd3f5e5), .K10_C14_W3(32'h3d151a31), .K10_C14_W4(32'hbd92031f), .K10_C14_W5(32'h3d37c885), .K10_C14_W6(32'h3ddbd864), .K10_C14_W7(32'hbdd1c93f), .K10_C14_W8(32'h3c1370bb), 
		.K10_C15_W0(32'h3d1a525f), .K10_C15_W1(32'hbde05ed3), .K10_C15_W2(32'hbd21b73b), .K10_C15_W3(32'hbceab915), .K10_C15_W4(32'hbdedef92), .K10_C15_W5(32'hbcf12129), .K10_C15_W6(32'h3d3fc6fd), .K10_C15_W7(32'hbd28dc76), .K10_C15_W8(32'hbe221980), 
		.K10_BIAS (32'h3d56fde2),

		.K11_C0_W0(32'hbdd79ee6), .K11_C0_W1(32'hbd73fee2), .K11_C0_W2(32'h3c80430b), .K11_C0_W3(32'h3cdff971), .K11_C0_W4(32'hbd9aaf4b), .K11_C0_W5(32'hbd0b35dc), .K11_C0_W6(32'hbddd88c1), .K11_C0_W7(32'h3df6f2a8), .K11_C0_W8(32'h3d92cf97), 
		.K11_C1_W0(32'h3e248ad8), .K11_C1_W1(32'hbddb0fde), .K11_C1_W2(32'h3cdfbb8c), .K11_C1_W3(32'h3cd86146), .K11_C1_W4(32'h3e043630), .K11_C1_W5(32'hbcecc97c), .K11_C1_W6(32'hbd4d91a6), .K11_C1_W7(32'hbd655def), .K11_C1_W8(32'hbe02ecbc), 
		.K11_C2_W0(32'hbdc02eab), .K11_C2_W1(32'h3e041ebe), .K11_C2_W2(32'h3d4917c5), .K11_C2_W3(32'h3e05a51f), .K11_C2_W4(32'h3cb66c05), .K11_C2_W5(32'h3d5b04db), .K11_C2_W6(32'hbdead507), .K11_C2_W7(32'h3db23f62), .K11_C2_W8(32'hbd90549d), 
		.K11_C3_W0(32'h3da058e4), .K11_C3_W1(32'h3e1ea787), .K11_C3_W2(32'h3d912e82), .K11_C3_W3(32'hbcb55572), .K11_C3_W4(32'hbe31e2d4), .K11_C3_W5(32'hbe128197), .K11_C3_W6(32'hbd2b8ed1), .K11_C3_W7(32'h3b0d0de6), .K11_C3_W8(32'hbcbc805d), 
		.K11_C4_W0(32'hbd3d31a8), .K11_C4_W1(32'h3c30e172), .K11_C4_W2(32'hbda70195), .K11_C4_W3(32'h3d366abd), .K11_C4_W4(32'h3dd89850), .K11_C4_W5(32'h3df255cd), .K11_C4_W6(32'hbca51794), .K11_C4_W7(32'h3e0786ae), .K11_C4_W8(32'h3afe3ddb), 
		.K11_C5_W0(32'hbdf3cde4), .K11_C5_W1(32'h3de5a6fc), .K11_C5_W2(32'h3c9900aa), .K11_C5_W3(32'h3d9776b8), .K11_C5_W4(32'h3e2e480b), .K11_C5_W5(32'h3e0b2219), .K11_C5_W6(32'h3e3164a3), .K11_C5_W7(32'h3db2d1ec), .K11_C5_W8(32'h3d90d7c6), 
		.K11_C6_W0(32'hbd86813f), .K11_C6_W1(32'hbd77022b), .K11_C6_W2(32'hbc8af92f), .K11_C6_W3(32'h3d741139), .K11_C6_W4(32'hbdbf719b), .K11_C6_W5(32'hbd7a8700), .K11_C6_W6(32'h3d1b5e47), .K11_C6_W7(32'hbd53fed1), .K11_C6_W8(32'hbdd637be), 
		.K11_C7_W0(32'h3db64db7), .K11_C7_W1(32'h3c5e153b), .K11_C7_W2(32'h3e014bcd), .K11_C7_W3(32'hbb5072d7), .K11_C7_W4(32'h3e1bfd80), .K11_C7_W5(32'hbd7ab3a9), .K11_C7_W6(32'hbd124941), .K11_C7_W7(32'hbcd1b9ad), .K11_C7_W8(32'h3e0c2b7b), 
		.K11_C8_W0(32'h3d2ab8f2), .K11_C8_W1(32'hbe20e20c), .K11_C8_W2(32'hbcfb7196), .K11_C8_W3(32'h3d5eb172), .K11_C8_W4(32'hbd165493), .K11_C8_W5(32'hbe45cec0), .K11_C8_W6(32'h3d92a768), .K11_C8_W7(32'hbd74c509), .K11_C8_W8(32'hbe1dda36), 
		.K11_C9_W0(32'h3c7a0bc7), .K11_C9_W1(32'h3d852e82), .K11_C9_W2(32'h3dd73707), .K11_C9_W3(32'h3e2e895a), .K11_C9_W4(32'h3e314c07), .K11_C9_W5(32'h3d90f9fa), .K11_C9_W6(32'h3dbcfe90), .K11_C9_W7(32'h3e021441), .K11_C9_W8(32'hbda0f6d1), 
		.K11_C10_W0(32'h3c6f27a1), .K11_C10_W1(32'hbd1c3ebf), .K11_C10_W2(32'h3dd424ff), .K11_C10_W3(32'h3dba32f7), .K11_C10_W4(32'hbda65ce5), .K11_C10_W5(32'h3e27b9cd), .K11_C10_W6(32'hbe1df3f3), .K11_C10_W7(32'h3e09afd8), .K11_C10_W8(32'h3d02eaf9), 
		.K11_C11_W0(32'hbe1d06f3), .K11_C11_W1(32'h3d399690), .K11_C11_W2(32'h3d0d5408), .K11_C11_W3(32'hbe0e4c68), .K11_C11_W4(32'h3d084219), .K11_C11_W5(32'hbd3b9d67), .K11_C11_W6(32'hbd0f4a68), .K11_C11_W7(32'hbc82ab63), .K11_C11_W8(32'h3dada66c), 
		.K11_C12_W0(32'h3dab916f), .K11_C12_W1(32'h3d4754a3), .K11_C12_W2(32'h3d19c190), .K11_C12_W3(32'h3e1d5dae), .K11_C12_W4(32'hbc711eff), .K11_C12_W5(32'h3e0ed7e8), .K11_C12_W6(32'h3e16bf29), .K11_C12_W7(32'hbdc99859), .K11_C12_W8(32'h3de7ba1d), 
		.K11_C13_W0(32'hbdf4454d), .K11_C13_W1(32'h3d9affd3), .K11_C13_W2(32'h3e09ce87), .K11_C13_W3(32'hbc9d09cf), .K11_C13_W4(32'hbd5b62eb), .K11_C13_W5(32'hbd22ad9f), .K11_C13_W6(32'hbd45b118), .K11_C13_W7(32'h3dcd7cd9), .K11_C13_W8(32'hbd7a28c8), 
		.K11_C14_W0(32'h3dbbe5eb), .K11_C14_W1(32'h3c8f17ff), .K11_C14_W2(32'hbd951054), .K11_C14_W3(32'h3c341025), .K11_C14_W4(32'hbda44e3b), .K11_C14_W5(32'h3d97d640), .K11_C14_W6(32'h3de259d9), .K11_C14_W7(32'hbda212a4), .K11_C14_W8(32'hbd57841d), 
		.K11_C15_W0(32'hbc9df2a1), .K11_C15_W1(32'hbdc6861a), .K11_C15_W2(32'hbe15a8a1), .K11_C15_W3(32'hbd9b790f), .K11_C15_W4(32'hbc325b3a), .K11_C15_W5(32'hbbddfb92), .K11_C15_W6(32'h3ddd4d7b), .K11_C15_W7(32'h3dec38c3), .K11_C15_W8(32'h3de37d00), 
		.K11_BIAS (32'hbc77a5c7),

		.K12_C0_W0(32'hbceb671d), .K12_C0_W1(32'hbd17e04b), .K12_C0_W2(32'hbdab3965), .K12_C0_W3(32'h3d3c09ca), .K12_C0_W4(32'h3c462efb), .K12_C0_W5(32'hbd4f7e32), .K12_C0_W6(32'h3de5c30c), .K12_C0_W7(32'h3d9d68a9), .K12_C0_W8(32'hbd7b3b9a), 
		.K12_C1_W0(32'hbdbf9ff3), .K12_C1_W1(32'hbd1fced6), .K12_C1_W2(32'h3da9db84), .K12_C1_W3(32'hbdca713d), .K12_C1_W4(32'h3dde71b1), .K12_C1_W5(32'hbbf72e1a), .K12_C1_W6(32'h3dd4f1c3), .K12_C1_W7(32'hbd90cf66), .K12_C1_W8(32'h3d9812c8), 
		.K12_C2_W0(32'hbc17eb5e), .K12_C2_W1(32'hbd84940f), .K12_C2_W2(32'hbd067f47), .K12_C2_W3(32'hbd7e78df), .K12_C2_W4(32'hbc9ff4ba), .K12_C2_W5(32'hbc4d3211), .K12_C2_W6(32'h3d776d04), .K12_C2_W7(32'hbe2cebd3), .K12_C2_W8(32'h3cf3206e), 
		.K12_C3_W0(32'hbc6f1035), .K12_C3_W1(32'h3cde338b), .K12_C3_W2(32'h3dd10c4b), .K12_C3_W3(32'hbd83c1ba), .K12_C3_W4(32'hbe207065), .K12_C3_W5(32'hbdaa05c7), .K12_C3_W6(32'h3d70b9dd), .K12_C3_W7(32'h3cae9d3d), .K12_C3_W8(32'hbdee5139), 
		.K12_C4_W0(32'hbe008256), .K12_C4_W1(32'hbc8eff7e), .K12_C4_W2(32'hbdb20df7), .K12_C4_W3(32'hbcc95080), .K12_C4_W4(32'hbdbe7713), .K12_C4_W5(32'h3df438eb), .K12_C4_W6(32'h3dd6538d), .K12_C4_W7(32'hbc8ed497), .K12_C4_W8(32'hbd5478ac), 
		.K12_C5_W0(32'hbd8d6c5f), .K12_C5_W1(32'h3dfcfc32), .K12_C5_W2(32'hbd6213a6), .K12_C5_W3(32'h3da54fb1), .K12_C5_W4(32'h3e0d23ee), .K12_C5_W5(32'h3e1b797b), .K12_C5_W6(32'h3e2bf9f9), .K12_C5_W7(32'hbdf2a124), .K12_C5_W8(32'h3d88bbc5), 
		.K12_C6_W0(32'hbe04fbb8), .K12_C6_W1(32'h3d617d52), .K12_C6_W2(32'hbd805094), .K12_C6_W3(32'h3dbae349), .K12_C6_W4(32'h3dbb549a), .K12_C6_W5(32'hbd3d3f39), .K12_C6_W6(32'h3e227298), .K12_C6_W7(32'h3dcd9cbe), .K12_C6_W8(32'h3d8bad63), 
		.K12_C7_W0(32'hbc8be555), .K12_C7_W1(32'h3ddbcfa7), .K12_C7_W2(32'h3d0d9fd7), .K12_C7_W3(32'h3db17fea), .K12_C7_W4(32'h3d4be78d), .K12_C7_W5(32'h3a99fd1f), .K12_C7_W6(32'hbbf1d53a), .K12_C7_W7(32'hbd93d5d6), .K12_C7_W8(32'hbc85ef12), 
		.K12_C8_W0(32'hbd7c0cc9), .K12_C8_W1(32'hbd427d83), .K12_C8_W2(32'h3d26acb9), .K12_C8_W3(32'h3ce8a4ca), .K12_C8_W4(32'h3c7be38f), .K12_C8_W5(32'h3c95776b), .K12_C8_W6(32'hbc5dcd53), .K12_C8_W7(32'h3d1b1c1d), .K12_C8_W8(32'hbc98376e), 
		.K12_C9_W0(32'h3dd4126c), .K12_C9_W1(32'h3de9a499), .K12_C9_W2(32'h3e030dee), .K12_C9_W3(32'hbd985489), .K12_C9_W4(32'h3e40da31), .K12_C9_W5(32'hbd47de90), .K12_C9_W6(32'h3d95a4a8), .K12_C9_W7(32'hbd562bbe), .K12_C9_W8(32'h3da79e01), 
		.K12_C10_W0(32'h3c5b3e0e), .K12_C10_W1(32'h3dad5af1), .K12_C10_W2(32'h3e1a2890), .K12_C10_W3(32'h3d8388e7), .K12_C10_W4(32'h3dffdb5c), .K12_C10_W5(32'hbd9d55e3), .K12_C10_W6(32'h3d74ee70), .K12_C10_W7(32'hbe05bbcb), .K12_C10_W8(32'hbcf0dfbd), 
		.K12_C11_W0(32'hbdc6fb42), .K12_C11_W1(32'h3c8d9d6a), .K12_C11_W2(32'h3e13a317), .K12_C11_W3(32'hbc0db81e), .K12_C11_W4(32'h3d283b43), .K12_C11_W5(32'hbd97c1e8), .K12_C11_W6(32'hbd4a3aa4), .K12_C11_W7(32'h3c0ef71f), .K12_C11_W8(32'h3dff8202), 
		.K12_C12_W0(32'h3dc78cd8), .K12_C12_W1(32'h3dd4afc7), .K12_C12_W2(32'h3d2edad7), .K12_C12_W3(32'hbddf18ad), .K12_C12_W4(32'h3d65d6fd), .K12_C12_W5(32'h3d190b8a), .K12_C12_W6(32'hbde0510e), .K12_C12_W7(32'hbe06b6d8), .K12_C12_W8(32'h3deeb1fe), 
		.K12_C13_W0(32'hbdd675d7), .K12_C13_W1(32'hbe10a2f7), .K12_C13_W2(32'h3d9a6af4), .K12_C13_W3(32'hbdc082a8), .K12_C13_W4(32'h3d20500b), .K12_C13_W5(32'hbd6af25d), .K12_C13_W6(32'h3d82a9e2), .K12_C13_W7(32'hbe0355e0), .K12_C13_W8(32'h3ddf93a8), 
		.K12_C14_W0(32'hbd892b72), .K12_C14_W1(32'h3e02ec85), .K12_C14_W2(32'h3dbc25c5), .K12_C14_W3(32'h3dbad981), .K12_C14_W4(32'hbe0c332f), .K12_C14_W5(32'hbdfff891), .K12_C14_W6(32'hbda1155a), .K12_C14_W7(32'h3e013d10), .K12_C14_W8(32'hbda158e7), 
		.K12_C15_W0(32'hbd0b1609), .K12_C15_W1(32'hbdf37951), .K12_C15_W2(32'hbe172fa3), .K12_C15_W3(32'h3d80830f), .K12_C15_W4(32'h3e15c4dc), .K12_C15_W5(32'hbb98d4c5), .K12_C15_W6(32'h3dbe1e59), .K12_C15_W7(32'hbdbb9c21), .K12_C15_W8(32'h3dfc5432), 
		.K12_BIAS (32'hbc8106b6),

		.K13_C0_W0(32'hbe01aaec), .K13_C0_W1(32'h3db4dbf6), .K13_C0_W2(32'hbca1931f), .K13_C0_W3(32'h3d1c9413), .K13_C0_W4(32'hbde8087e), .K13_C0_W5(32'hbd8bfcaf), .K13_C0_W6(32'h3e006631), .K13_C0_W7(32'hbe009a6a), .K13_C0_W8(32'hbc2538e2), 
		.K13_C1_W0(32'hbdb97fab), .K13_C1_W1(32'h3cc1cda4), .K13_C1_W2(32'h3c244d1f), .K13_C1_W3(32'h3d839ffe), .K13_C1_W4(32'hbd9d8ba4), .K13_C1_W5(32'hbbb9d666), .K13_C1_W6(32'h3c5a615e), .K13_C1_W7(32'h3c983408), .K13_C1_W8(32'hbe04980e), 
		.K13_C2_W0(32'h3dacf76d), .K13_C2_W1(32'hbe04bb09), .K13_C2_W2(32'hbd01986d), .K13_C2_W3(32'hbdefd094), .K13_C2_W4(32'hbbc59c6f), .K13_C2_W5(32'h3dd4e0ee), .K13_C2_W6(32'h3df55aed), .K13_C2_W7(32'h3d48d74e), .K13_C2_W8(32'hbe00fe71), 
		.K13_C3_W0(32'hbcb05513), .K13_C3_W1(32'h3d019709), .K13_C3_W2(32'h3c22bbd0), .K13_C3_W3(32'h3ccfca09), .K13_C3_W4(32'hbcda8630), .K13_C3_W5(32'hbde84cfc), .K13_C3_W6(32'hbdfbd6e3), .K13_C3_W7(32'h3d9ac6f4), .K13_C3_W8(32'hbda31bb1), 
		.K13_C4_W0(32'h3d480de7), .K13_C4_W1(32'hbcdae26e), .K13_C4_W2(32'hbcf9c658), .K13_C4_W3(32'h3d928cc9), .K13_C4_W4(32'h3df55988), .K13_C4_W5(32'h3d6f1d04), .K13_C4_W6(32'h3db4d8fd), .K13_C4_W7(32'h3c13af34), .K13_C4_W8(32'hbb49cb67), 
		.K13_C5_W0(32'h3e3b1a03), .K13_C5_W1(32'hbab50904), .K13_C5_W2(32'h3df66bf3), .K13_C5_W3(32'hbdff6273), .K13_C5_W4(32'h3d133daf), .K13_C5_W5(32'h3d8aba51), .K13_C5_W6(32'hbc7e3dd9), .K13_C5_W7(32'h3dc020b2), .K13_C5_W8(32'hbd78cf13), 
		.K13_C6_W0(32'hbce9ebd6), .K13_C6_W1(32'h3db83730), .K13_C6_W2(32'hbdbf8058), .K13_C6_W3(32'h3e10d1a5), .K13_C6_W4(32'hbe0d354b), .K13_C6_W5(32'h3c8090ea), .K13_C6_W6(32'hbcb2355e), .K13_C6_W7(32'h3c11d9a5), .K13_C6_W8(32'hbe17c7a1), 
		.K13_C7_W0(32'h3da516bd), .K13_C7_W1(32'hbc15098e), .K13_C7_W2(32'hbe0acde6), .K13_C7_W3(32'hbbe1347a), .K13_C7_W4(32'h3dc67ec1), .K13_C7_W5(32'h3d059603), .K13_C7_W6(32'hbddc25e6), .K13_C7_W7(32'h3b437d90), .K13_C7_W8(32'h3da284a4), 
		.K13_C8_W0(32'h3dc911a8), .K13_C8_W1(32'hbe21f9ea), .K13_C8_W2(32'h3d56b6f3), .K13_C8_W3(32'h3c72af11), .K13_C8_W4(32'hbde19b27), .K13_C8_W5(32'hbcc3b95e), .K13_C8_W6(32'hbcb399f1), .K13_C8_W7(32'h3dd39d6c), .K13_C8_W8(32'hbdb53799), 
		.K13_C9_W0(32'h3cd8e57b), .K13_C9_W1(32'h3e3872a4), .K13_C9_W2(32'h3ded5aae), .K13_C9_W3(32'h3db50300), .K13_C9_W4(32'hbdf6dbfe), .K13_C9_W5(32'h3de50d1f), .K13_C9_W6(32'h3db5f4eb), .K13_C9_W7(32'h3ca9e8b6), .K13_C9_W8(32'hbd6b2adc), 
		.K13_C10_W0(32'h3caa2978), .K13_C10_W1(32'h3bf25353), .K13_C10_W2(32'h3df85293), .K13_C10_W3(32'h3d00bfbf), .K13_C10_W4(32'h3d861e4c), .K13_C10_W5(32'h3de5cfab), .K13_C10_W6(32'hbd9e828a), .K13_C10_W7(32'hbdea50c2), .K13_C10_W8(32'h3da4ff79), 
		.K13_C11_W0(32'h3d6db93f), .K13_C11_W1(32'h3dd0360f), .K13_C11_W2(32'hbc1ecedf), .K13_C11_W3(32'h3dcd50e5), .K13_C11_W4(32'hbe00db58), .K13_C11_W5(32'hbd086ee3), .K13_C11_W6(32'hbd8fa079), .K13_C11_W7(32'h3d8e1f43), .K13_C11_W8(32'hbd7287bb), 
		.K13_C12_W0(32'hbdb20654), .K13_C12_W1(32'h3d6c53d7), .K13_C12_W2(32'h3dc4df3c), .K13_C12_W3(32'h3e2361b7), .K13_C12_W4(32'h3dd22d62), .K13_C12_W5(32'hbdc6782d), .K13_C12_W6(32'h3d6c5f11), .K13_C12_W7(32'hbd75fd72), .K13_C12_W8(32'hbd8ae985), 
		.K13_C13_W0(32'hbdecb627), .K13_C13_W1(32'hbd88245b), .K13_C13_W2(32'h3debd99f), .K13_C13_W3(32'hbdda2eb2), .K13_C13_W4(32'hbdf2d93a), .K13_C13_W5(32'h3dd056ed), .K13_C13_W6(32'h3d365823), .K13_C13_W7(32'h3de4d5f3), .K13_C13_W8(32'h3dc14af5), 
		.K13_C14_W0(32'h3dacffeb), .K13_C14_W1(32'hbe03704b), .K13_C14_W2(32'h3d69c7f9), .K13_C14_W3(32'h3aa809b8), .K13_C14_W4(32'hbda0842e), .K13_C14_W5(32'h3db39afa), .K13_C14_W6(32'h3d9f3c4f), .K13_C14_W7(32'hbcc66ca4), .K13_C14_W8(32'h39569f5f), 
		.K13_C15_W0(32'h3de5f5ba), .K13_C15_W1(32'h3c90a6fe), .K13_C15_W2(32'hbdfced58), .K13_C15_W3(32'h3df7e9b2), .K13_C15_W4(32'h3d11bb75), .K13_C15_W5(32'h3d7b96de), .K13_C15_W6(32'hbb575a56), .K13_C15_W7(32'hbd220491), .K13_C15_W8(32'hbc44fcb2), 
		.K13_BIAS (32'hbbc561ac),

		.K14_C0_W0(32'h3e015c2d), .K14_C0_W1(32'hbab7df3b), .K14_C0_W2(32'h3d494539), .K14_C0_W3(32'h3dae0a61), .K14_C0_W4(32'h3de8e85a), .K14_C0_W5(32'h3d9be73e), .K14_C0_W6(32'h3df5156b), .K14_C0_W7(32'hbc67a204), .K14_C0_W8(32'h3d4edc13), 
		.K14_C1_W0(32'hbdf864b1), .K14_C1_W1(32'h3d1a6880), .K14_C1_W2(32'hbdf55c16), .K14_C1_W3(32'hbdf49616), .K14_C1_W4(32'hbe1173fd), .K14_C1_W5(32'h3dfacf24), .K14_C1_W6(32'hbe0c4d22), .K14_C1_W7(32'h3cf7b88e), .K14_C1_W8(32'h3bdaf1f9), 
		.K14_C2_W0(32'hbdf431d3), .K14_C2_W1(32'hbde4b14d), .K14_C2_W2(32'h3e082dd5), .K14_C2_W3(32'hbd4c6721), .K14_C2_W4(32'h3d7df34f), .K14_C2_W5(32'hbdf47991), .K14_C2_W6(32'h3d8d256e), .K14_C2_W7(32'h3d77f5a9), .K14_C2_W8(32'h3da33e25), 
		.K14_C3_W0(32'h3e1792fd), .K14_C3_W1(32'h3e09564b), .K14_C3_W2(32'h3d4a5ac9), .K14_C3_W3(32'h3ce4f3a6), .K14_C3_W4(32'hbd897cfc), .K14_C3_W5(32'hbe020767), .K14_C3_W6(32'h3d49e3eb), .K14_C3_W7(32'h3d4ff6d3), .K14_C3_W8(32'hbd18da19), 
		.K14_C4_W0(32'h3d7eaf6a), .K14_C4_W1(32'hbdeb6a4d), .K14_C4_W2(32'h3def3617), .K14_C4_W3(32'hbdb71748), .K14_C4_W4(32'hbdd5e467), .K14_C4_W5(32'hbdc8c21d), .K14_C4_W6(32'hbe1a8427), .K14_C4_W7(32'hbdfcb9f7), .K14_C4_W8(32'hbe097c88), 
		.K14_C5_W0(32'hbde8d460), .K14_C5_W1(32'hbd429987), .K14_C5_W2(32'hbd6d05a6), .K14_C5_W3(32'hbae5292d), .K14_C5_W4(32'hbde49b40), .K14_C5_W5(32'h3ce520f4), .K14_C5_W6(32'hbe082d1b), .K14_C5_W7(32'h3dbc7e5d), .K14_C5_W8(32'h3dab9361), 
		.K14_C6_W0(32'hbd2ab6f0), .K14_C6_W1(32'h3d928ce2), .K14_C6_W2(32'h3d9655c2), .K14_C6_W3(32'h3d173e0a), .K14_C6_W4(32'hbd8e3708), .K14_C6_W5(32'h3db18c60), .K14_C6_W6(32'hbc05f58a), .K14_C6_W7(32'hbdc390ab), .K14_C6_W8(32'hbdb05a76), 
		.K14_C7_W0(32'hbdec3a33), .K14_C7_W1(32'h3d925b6e), .K14_C7_W2(32'h3c5c32f1), .K14_C7_W3(32'hbd998d75), .K14_C7_W4(32'h3e071be2), .K14_C7_W5(32'hbd269853), .K14_C7_W6(32'hbdfb68f3), .K14_C7_W7(32'hbc427542), .K14_C7_W8(32'h3cc588a8), 
		.K14_C8_W0(32'hbd990860), .K14_C8_W1(32'hbdc76524), .K14_C8_W2(32'hbd223247), .K14_C8_W3(32'h3db57da7), .K14_C8_W4(32'h3da4fb07), .K14_C8_W5(32'h3e0feadd), .K14_C8_W6(32'h3e10644a), .K14_C8_W7(32'h3d2ca52d), .K14_C8_W8(32'hbe091196), 
		.K14_C9_W0(32'h3e076292), .K14_C9_W1(32'h3d10a3f4), .K14_C9_W2(32'h3d3e22ce), .K14_C9_W3(32'h3e07b3e1), .K14_C9_W4(32'hbc8589d3), .K14_C9_W5(32'hbdd9062f), .K14_C9_W6(32'h3cfa7086), .K14_C9_W7(32'h3d9d05c3), .K14_C9_W8(32'hbdd2f8e2), 
		.K14_C10_W0(32'h3c994966), .K14_C10_W1(32'hbdcf07c2), .K14_C10_W2(32'h3d6e9cb8), .K14_C10_W3(32'hbddb75fc), .K14_C10_W4(32'h3e05fec6), .K14_C10_W5(32'h3c05becc), .K14_C10_W6(32'hbde1128a), .K14_C10_W7(32'h3d57cadc), .K14_C10_W8(32'hbe0800dc), 
		.K14_C11_W0(32'h3dd8e42f), .K14_C11_W1(32'hbdb71625), .K14_C11_W2(32'hbd92b5b9), .K14_C11_W3(32'hbdc21d56), .K14_C11_W4(32'hbdaa05d0), .K14_C11_W5(32'hbd388dde), .K14_C11_W6(32'h3e262014), .K14_C11_W7(32'h3dc05524), .K14_C11_W8(32'hbde57cb5), 
		.K14_C12_W0(32'h3db92a58), .K14_C12_W1(32'hbdbda618), .K14_C12_W2(32'hbd17e909), .K14_C12_W3(32'h3d047afb), .K14_C12_W4(32'h3db15524), .K14_C12_W5(32'h3e00d644), .K14_C12_W6(32'hbdcf09b5), .K14_C12_W7(32'h3d8c2b29), .K14_C12_W8(32'hbc78e5f6), 
		.K14_C13_W0(32'h3b0dc631), .K14_C13_W1(32'hbd9f9a6d), .K14_C13_W2(32'hbd6c7f0c), .K14_C13_W3(32'h3df17358), .K14_C13_W4(32'hbd4cba02), .K14_C13_W5(32'h3e00fa46), .K14_C13_W6(32'hbe15ca22), .K14_C13_W7(32'hbd7921e9), .K14_C13_W8(32'h3c9596d5), 
		.K14_C14_W0(32'hbd9789b6), .K14_C14_W1(32'hbbe74655), .K14_C14_W2(32'h3d9c6a9e), .K14_C14_W3(32'hbdc2597d), .K14_C14_W4(32'hbd77a926), .K14_C14_W5(32'h3d642846), .K14_C14_W6(32'h3dbe9520), .K14_C14_W7(32'h3d126987), .K14_C14_W8(32'h3d6d34da), 
		.K14_C15_W0(32'hbd656154), .K14_C15_W1(32'hbd443775), .K14_C15_W2(32'hbdfd9ad5), .K14_C15_W3(32'h3d52919c), .K14_C15_W4(32'h3d4f956d), .K14_C15_W5(32'hbca34dc4), .K14_C15_W6(32'hbdd2d077), .K14_C15_W7(32'h3dfc9f0f), .K14_C15_W8(32'hbdc42bf7), 
		.K14_BIAS (32'hba8b09b8),

		.K15_C0_W0(32'h3d592cb4), .K15_C0_W1(32'h3db45944), .K15_C0_W2(32'h3c94ae72), .K15_C0_W3(32'hbe0f1aa8), .K15_C0_W4(32'hbc120a59), .K15_C0_W5(32'h3de49053), .K15_C0_W6(32'hbdf4e055), .K15_C0_W7(32'hbc9d1fff), .K15_C0_W8(32'h3b007f27), 
		.K15_C1_W0(32'hbdc1fb66), .K15_C1_W1(32'h3db91141), .K15_C1_W2(32'h3dfcd166), .K15_C1_W3(32'hbb2205cf), .K15_C1_W4(32'hbe1eb115), .K15_C1_W5(32'hb95fed70), .K15_C1_W6(32'hbca9e780), .K15_C1_W7(32'hba75e614), .K15_C1_W8(32'h3e0ecf46), 
		.K15_C2_W0(32'hbdf69809), .K15_C2_W1(32'hbd28d3fe), .K15_C2_W2(32'hbe1842b5), .K15_C2_W3(32'hbd99fadf), .K15_C2_W4(32'hbd0ff8e5), .K15_C2_W5(32'h3e003eff), .K15_C2_W6(32'hbc4bbb0a), .K15_C2_W7(32'h3d9eeaf2), .K15_C2_W8(32'hbc02dfe6), 
		.K15_C3_W0(32'h3d077783), .K15_C3_W1(32'h3cbd2aa4), .K15_C3_W2(32'hbe1c3217), .K15_C3_W3(32'hbd8076d8), .K15_C3_W4(32'hbd70417f), .K15_C3_W5(32'h3d230160), .K15_C3_W6(32'hbdc1bc84), .K15_C3_W7(32'h3bd43585), .K15_C3_W8(32'hbdb090fc), 
		.K15_C4_W0(32'hbd2a445e), .K15_C4_W1(32'h3d9d6a7c), .K15_C4_W2(32'hbd9cec9e), .K15_C4_W3(32'h3cd50a83), .K15_C4_W4(32'h3d40762b), .K15_C4_W5(32'h3d62fa1f), .K15_C4_W6(32'h3da432fd), .K15_C4_W7(32'h3da9fd26), .K15_C4_W8(32'h3d5b108e), 
		.K15_C5_W0(32'h3db5473e), .K15_C5_W1(32'h3e191e41), .K15_C5_W2(32'hbdea2953), .K15_C5_W3(32'h3e100ce2), .K15_C5_W4(32'h3df6eab1), .K15_C5_W5(32'hbd8692d7), .K15_C5_W6(32'h3df153d4), .K15_C5_W7(32'h3dbd3b54), .K15_C5_W8(32'hbdc3903d), 
		.K15_C6_W0(32'hbe442341), .K15_C6_W1(32'hbdebd043), .K15_C6_W2(32'hbc931733), .K15_C6_W3(32'h3d0f97ec), .K15_C6_W4(32'hbd5eb56f), .K15_C6_W5(32'h3d87f4b1), .K15_C6_W6(32'hbd4c3bef), .K15_C6_W7(32'hbdb00b68), .K15_C6_W8(32'hbc828f87), 
		.K15_C7_W0(32'hbdccd572), .K15_C7_W1(32'h3d36ecf8), .K15_C7_W2(32'hbdad168e), .K15_C7_W3(32'hbdd6743d), .K15_C7_W4(32'h3e013c34), .K15_C7_W5(32'hbdd7faad), .K15_C7_W6(32'hbdce3701), .K15_C7_W7(32'h3b81186e), .K15_C7_W8(32'h3d2423a8), 
		.K15_C8_W0(32'h3d9d69cd), .K15_C8_W1(32'h3df33603), .K15_C8_W2(32'hbd6d8bed), .K15_C8_W3(32'h3e28816a), .K15_C8_W4(32'hbdfed1ae), .K15_C8_W5(32'h3e07de63), .K15_C8_W6(32'h3d6bf2c2), .K15_C8_W7(32'h3df13380), .K15_C8_W8(32'h3e09e091), 
		.K15_C9_W0(32'h3c60d546), .K15_C9_W1(32'hbe023e61), .K15_C9_W2(32'h3d11fafc), .K15_C9_W3(32'h3d9cf61c), .K15_C9_W4(32'h3d44fcbf), .K15_C9_W5(32'h3da77da8), .K15_C9_W6(32'h3d362d6e), .K15_C9_W7(32'h3de89e85), .K15_C9_W8(32'h3d9c7655), 
		.K15_C10_W0(32'hbde457b3), .K15_C10_W1(32'hbd9ecadb), .K15_C10_W2(32'h3d326ed0), .K15_C10_W3(32'h3d82ed66), .K15_C10_W4(32'hbdf9dcf4), .K15_C10_W5(32'h3d59fe3e), .K15_C10_W6(32'hbdc91ef8), .K15_C10_W7(32'hbb2d86cc), .K15_C10_W8(32'h3c978ac3), 
		.K15_C11_W0(32'hbdace967), .K15_C11_W1(32'hbdb8bd9b), .K15_C11_W2(32'h3d4067a8), .K15_C11_W3(32'hbdf5f43d), .K15_C11_W4(32'hbbae1912), .K15_C11_W5(32'h3d7032e5), .K15_C11_W6(32'h3e10d406), .K15_C11_W7(32'h3dbffacb), .K15_C11_W8(32'hbd941686), 
		.K15_C12_W0(32'h3d9206e8), .K15_C12_W1(32'hbd383df8), .K15_C12_W2(32'hbd32b00b), .K15_C12_W3(32'h3cfd01fe), .K15_C12_W4(32'hbdf87ae2), .K15_C12_W5(32'hbd670e56), .K15_C12_W6(32'h3daa780f), .K15_C12_W7(32'hbe017f94), .K15_C12_W8(32'h3d8aae76), 
		.K15_C13_W0(32'h3c8d03da), .K15_C13_W1(32'h3df647f4), .K15_C13_W2(32'h3deeedc0), .K15_C13_W3(32'hbdccdb58), .K15_C13_W4(32'h3ccf6b1a), .K15_C13_W5(32'h3df50af7), .K15_C13_W6(32'h3cfcb42e), .K15_C13_W7(32'hbd53911e), .K15_C13_W8(32'hbd4f3734), 
		.K15_C14_W0(32'h3e366cb8), .K15_C14_W1(32'h3e01a973), .K15_C14_W2(32'h3d053db6), .K15_C14_W3(32'h3e1389fe), .K15_C14_W4(32'hbd337b1d), .K15_C14_W5(32'hbdec5d87), .K15_C14_W6(32'hbdd6eccf), .K15_C14_W7(32'h3dd60c89), .K15_C14_W8(32'hbdfcbbe5), 
		.K15_C15_W0(32'h3e170e8f), .K15_C15_W1(32'hbdaaabb7), .K15_C15_W2(32'h3dd8b3db), .K15_C15_W3(32'hbdb1a0ae), .K15_C15_W4(32'h3ce9260b), .K15_C15_W5(32'hbdc46f69), .K15_C15_W6(32'hbdde7397), .K15_C15_W7(32'h3d9c14e1), .K15_C15_W8(32'hbdb93c15), 
		.K15_BIAS (32'h3d34f629)
		)
		block4_conv3(
		.clk(clk),
		.resetn(resetn),
		.data_valid_in(conv_valid_out_4_2),
		.data_in_0(conv_out_4_2[0]),
		.data_in_1(conv_out_4_2[1]),
		.data_in_2(conv_out_4_2[2]),
		.data_in_3(conv_out_4_2[3]),
		.data_in_4(conv_out_4_2[4]),
		.data_in_5(conv_out_4_2[5]),
		.data_in_6(conv_out_4_2[6]),
		.data_in_7(conv_out_4_2[7]),
		.data_in_8(conv_out_4_2[8]),
		.data_in_9(conv_out_4_2[9]),
		.data_in_10(conv_out_4_2[10]),
		.data_in_11(conv_out_4_2[11]),
		.data_in_12(conv_out_4_2[12]),
		.data_in_13(conv_out_4_2[13]),
		.data_in_14(conv_out_4_2[14]),
		.data_in_15(conv_out_4_2[15]),
		.data_out_conv_0(conv_out_4_3[0]),
		.data_out_conv_1(conv_out_4_3[1]),
		.data_out_conv_2(conv_out_4_3[2]),
		.data_out_conv_3(conv_out_4_3[3]),
		.data_out_conv_4(conv_out_4_3[4]),
		.data_out_conv_5(conv_out_4_3[5]),
		.data_out_conv_6(conv_out_4_3[6]),
		.data_out_conv_7(conv_out_4_3[7]),
		.data_out_conv_8(conv_out_4_3[8]),
		.data_out_conv_9(conv_out_4_3[9]),
		.data_out_conv_10(conv_out_4_3[10]),
		.data_out_conv_11(conv_out_4_3[11]),
		.data_out_conv_12(conv_out_4_3[12]),
		.data_out_conv_13(conv_out_4_3[13]),
		.data_out_conv_14(conv_out_4_3[14]),
		.data_out_conv_15(conv_out_4_3[15]),
		.valid_out_pixel(conv_valid_out_4_3),
		.done(done_conv_4_3)
		);



    genvar i;

    generate
    for (i = 0; i < CHANNEL_OUT; i=i+1) 
    begin : gen_relu // needs CHANNEL_OUT relu

        activate #(
            .DATA_WIDTH(32)
        )
        relu (
            .in(conv_out_4_3[i]),			// Edit here
            .out(relu_out[i])
        );
    end
    endgenerate

    generate
    for (i = 0; i < CHANNEL_OUT; i=i+1) 
    begin : gen_max_pool // needs CHANNEL_OUT max_pooling

        max_pooling #(
            .DATA_WIDTH(32),
            .WIDTH(WIDTH),
            .HEIGHT(HEIGHT)
        )
        max_pool(
            .clk(clk),
			.ack(done_conv_4_3),					// Edit here
            .resetn(resetn),
            .valid_in(conv_valid_out_4_3),			// Edit here
            .data_in(relu_out[i]),
            .data_out(data_out_pool[i]),
            .valid_out(valid_out_pool[i]),
            .done(done_pool[i])
        );
    end
    endgenerate

endmodule